`timescale 1ns / 1ps

module out_fifo_args (
    input acc_clk,
    input dm_clk,
    //control interface
    input aresetn,
    input out_fifo_allow,
    output [C_NUM_OUTPUT_FIFOs-1:0] out_fifo_ready,
    output [C_NUM_OUTPUT_FIFOs-1:0] out_fifo_finished,
    //output FIFO to AXI-Stream interface 0
    output m_axis_fifo_0_tlast,
    output m_axis_fifo_0_tvalid,
    output [C_OUTPUT_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tkeep,
    output [C_OUTPUT_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tstrb,
    output [C_OUTPUT_FIFO_0_DMWIDTH-1:0] m_axis_fifo_0_tdata,
    input m_axis_fifo_0_tready,
    output ap_fifo_oarg_0_full_n,
    input [C_OUTPUT_FIFO_0_WIDTH-1:0] ap_fifo_oarg_0_din,
    input ap_fifo_oarg_0_write,
    //output FIFO to AXI-Stream interface 1
    output m_axis_fifo_1_tlast,
    output m_axis_fifo_1_tvalid,
    output [C_OUTPUT_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tkeep,
    output [C_OUTPUT_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tstrb,
    output [C_OUTPUT_FIFO_1_DMWIDTH-1:0] m_axis_fifo_1_tdata,
    input m_axis_fifo_1_tready,
    output ap_fifo_oarg_1_full_n,
    input [C_OUTPUT_FIFO_1_WIDTH-1:0] ap_fifo_oarg_1_din,
    input ap_fifo_oarg_1_write,
    //output FIFO to AXI-Stream interface 2
    output m_axis_fifo_2_tlast,
    output m_axis_fifo_2_tvalid,
    output [C_OUTPUT_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tkeep,
    output [C_OUTPUT_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tstrb,
    output [C_OUTPUT_FIFO_2_DMWIDTH-1:0] m_axis_fifo_2_tdata,
    input m_axis_fifo_2_tready,
    output ap_fifo_oarg_2_full_n,
    input [C_OUTPUT_FIFO_2_WIDTH-1:0] ap_fifo_oarg_2_din,
    input ap_fifo_oarg_2_write,
    //output FIFO to AXI-Stream interface 3
    output m_axis_fifo_3_tlast,
    output m_axis_fifo_3_tvalid,
    output [C_OUTPUT_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tkeep,
    output [C_OUTPUT_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tstrb,
    output [C_OUTPUT_FIFO_3_DMWIDTH-1:0] m_axis_fifo_3_tdata,
    input m_axis_fifo_3_tready,
    output ap_fifo_oarg_3_full_n,
    input [C_OUTPUT_FIFO_3_WIDTH-1:0] ap_fifo_oarg_3_din,
    input ap_fifo_oarg_3_write,
    //output FIFO to AXI-Stream interface 4
    output m_axis_fifo_4_tlast,
    output m_axis_fifo_4_tvalid,
    output [C_OUTPUT_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tkeep,
    output [C_OUTPUT_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tstrb,
    output [C_OUTPUT_FIFO_4_DMWIDTH-1:0] m_axis_fifo_4_tdata,
    input m_axis_fifo_4_tready,
    output ap_fifo_oarg_4_full_n,
    input [C_OUTPUT_FIFO_4_WIDTH-1:0] ap_fifo_oarg_4_din,
    input ap_fifo_oarg_4_write,
    //output FIFO to AXI-Stream interface 5
    output m_axis_fifo_5_tlast,
    output m_axis_fifo_5_tvalid,
    output [C_OUTPUT_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tkeep,
    output [C_OUTPUT_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tstrb,
    output [C_OUTPUT_FIFO_5_DMWIDTH-1:0] m_axis_fifo_5_tdata,
    input m_axis_fifo_5_tready,
    output ap_fifo_oarg_5_full_n,
    input [C_OUTPUT_FIFO_5_WIDTH-1:0] ap_fifo_oarg_5_din,
    input ap_fifo_oarg_5_write,
    //output FIFO to AXI-Stream interface 6
    output m_axis_fifo_6_tlast,
    output m_axis_fifo_6_tvalid,
    output [C_OUTPUT_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tkeep,
    output [C_OUTPUT_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tstrb,
    output [C_OUTPUT_FIFO_6_DMWIDTH-1:0] m_axis_fifo_6_tdata,
    input m_axis_fifo_6_tready,
    output ap_fifo_oarg_6_full_n,
    input [C_OUTPUT_FIFO_6_WIDTH-1:0] ap_fifo_oarg_6_din,
    input ap_fifo_oarg_6_write,
    //output FIFO to AXI-Stream interface 7
    output m_axis_fifo_7_tlast,
    output m_axis_fifo_7_tvalid,
    output [C_OUTPUT_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tkeep,
    output [C_OUTPUT_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tstrb,
    output [C_OUTPUT_FIFO_7_DMWIDTH-1:0] m_axis_fifo_7_tdata,
    input m_axis_fifo_7_tready,
    output ap_fifo_oarg_7_full_n,
    input [C_OUTPUT_FIFO_7_WIDTH-1:0] ap_fifo_oarg_7_din,
    input ap_fifo_oarg_7_write,
    //output FIFO to AXI-Stream interface 8
    output m_axis_fifo_8_tlast,
    output m_axis_fifo_8_tvalid,
    output [C_OUTPUT_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tkeep,
    output [C_OUTPUT_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tstrb,
    output [C_OUTPUT_FIFO_8_DMWIDTH-1:0] m_axis_fifo_8_tdata,
    input m_axis_fifo_8_tready,
    output ap_fifo_oarg_8_full_n,
    input [C_OUTPUT_FIFO_8_WIDTH-1:0] ap_fifo_oarg_8_din,
    input ap_fifo_oarg_8_write,
    //output FIFO to AXI-Stream interface 9
    output m_axis_fifo_9_tlast,
    output m_axis_fifo_9_tvalid,
    output [C_OUTPUT_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tkeep,
    output [C_OUTPUT_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tstrb,
    output [C_OUTPUT_FIFO_9_DMWIDTH-1:0] m_axis_fifo_9_tdata,
    input m_axis_fifo_9_tready,
    output ap_fifo_oarg_9_full_n,
    input [C_OUTPUT_FIFO_9_WIDTH-1:0] ap_fifo_oarg_9_din,
    input ap_fifo_oarg_9_write,
    //output FIFO to AXI-Stream interface 10
    output m_axis_fifo_10_tlast,
    output m_axis_fifo_10_tvalid,
    output [C_OUTPUT_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tkeep,
    output [C_OUTPUT_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tstrb,
    output [C_OUTPUT_FIFO_10_DMWIDTH-1:0] m_axis_fifo_10_tdata,
    input m_axis_fifo_10_tready,
    output ap_fifo_oarg_10_full_n,
    input [C_OUTPUT_FIFO_10_WIDTH-1:0] ap_fifo_oarg_10_din,
    input ap_fifo_oarg_10_write,
    //output FIFO to AXI-Stream interface 11
    output m_axis_fifo_11_tlast,
    output m_axis_fifo_11_tvalid,
    output [C_OUTPUT_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tkeep,
    output [C_OUTPUT_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tstrb,
    output [C_OUTPUT_FIFO_11_DMWIDTH-1:0] m_axis_fifo_11_tdata,
    input m_axis_fifo_11_tready,
    output ap_fifo_oarg_11_full_n,
    input [C_OUTPUT_FIFO_11_WIDTH-1:0] ap_fifo_oarg_11_din,
    input ap_fifo_oarg_11_write,
    //output FIFO to AXI-Stream interface 12
    output m_axis_fifo_12_tlast,
    output m_axis_fifo_12_tvalid,
    output [C_OUTPUT_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tkeep,
    output [C_OUTPUT_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tstrb,
    output [C_OUTPUT_FIFO_12_DMWIDTH-1:0] m_axis_fifo_12_tdata,
    input m_axis_fifo_12_tready,
    output ap_fifo_oarg_12_full_n,
    input [C_OUTPUT_FIFO_12_WIDTH-1:0] ap_fifo_oarg_12_din,
    input ap_fifo_oarg_12_write,
    //output FIFO to AXI-Stream interface 13
    output m_axis_fifo_13_tlast,
    output m_axis_fifo_13_tvalid,
    output [C_OUTPUT_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tkeep,
    output [C_OUTPUT_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tstrb,
    output [C_OUTPUT_FIFO_13_DMWIDTH-1:0] m_axis_fifo_13_tdata,
    input m_axis_fifo_13_tready,
    output ap_fifo_oarg_13_full_n,
    input [C_OUTPUT_FIFO_13_WIDTH-1:0] ap_fifo_oarg_13_din,
    input ap_fifo_oarg_13_write,
    //output FIFO to AXI-Stream interface 14
    output m_axis_fifo_14_tlast,
    output m_axis_fifo_14_tvalid,
    output [C_OUTPUT_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tkeep,
    output [C_OUTPUT_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tstrb,
    output [C_OUTPUT_FIFO_14_DMWIDTH-1:0] m_axis_fifo_14_tdata,
    input m_axis_fifo_14_tready,
    output ap_fifo_oarg_14_full_n,
    input [C_OUTPUT_FIFO_14_WIDTH-1:0] ap_fifo_oarg_14_din,
    input ap_fifo_oarg_14_write,
    //output FIFO to AXI-Stream interface 15
    output m_axis_fifo_15_tlast,
    output m_axis_fifo_15_tvalid,
    output [C_OUTPUT_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tkeep,
    output [C_OUTPUT_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tstrb,
    output [C_OUTPUT_FIFO_15_DMWIDTH-1:0] m_axis_fifo_15_tdata,
    input m_axis_fifo_15_tready,
    output ap_fifo_oarg_15_full_n,
    input [C_OUTPUT_FIFO_15_WIDTH-1:0] ap_fifo_oarg_15_din,
    input ap_fifo_oarg_15_write,
    //output FIFO to AXI-Stream interface 16
    output m_axis_fifo_16_tlast,
    output m_axis_fifo_16_tvalid,
    output [C_OUTPUT_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tkeep,
    output [C_OUTPUT_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tstrb,
    output [C_OUTPUT_FIFO_16_DMWIDTH-1:0] m_axis_fifo_16_tdata,
    input m_axis_fifo_16_tready,
    output ap_fifo_oarg_16_full_n,
    input [C_OUTPUT_FIFO_16_WIDTH-1:0] ap_fifo_oarg_16_din,
    input ap_fifo_oarg_16_write,
    //output FIFO to AXI-Stream interface 17
    output m_axis_fifo_17_tlast,
    output m_axis_fifo_17_tvalid,
    output [C_OUTPUT_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tkeep,
    output [C_OUTPUT_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tstrb,
    output [C_OUTPUT_FIFO_17_DMWIDTH-1:0] m_axis_fifo_17_tdata,
    input m_axis_fifo_17_tready,
    output ap_fifo_oarg_17_full_n,
    input [C_OUTPUT_FIFO_17_WIDTH-1:0] ap_fifo_oarg_17_din,
    input ap_fifo_oarg_17_write,
    //output FIFO to AXI-Stream interface 18
    output m_axis_fifo_18_tlast,
    output m_axis_fifo_18_tvalid,
    output [C_OUTPUT_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tkeep,
    output [C_OUTPUT_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tstrb,
    output [C_OUTPUT_FIFO_18_DMWIDTH-1:0] m_axis_fifo_18_tdata,
    input m_axis_fifo_18_tready,
    output ap_fifo_oarg_18_full_n,
    input [C_OUTPUT_FIFO_18_WIDTH-1:0] ap_fifo_oarg_18_din,
    input ap_fifo_oarg_18_write,
    //output FIFO to AXI-Stream interface 19
    output m_axis_fifo_19_tlast,
    output m_axis_fifo_19_tvalid,
    output [C_OUTPUT_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tkeep,
    output [C_OUTPUT_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tstrb,
    output [C_OUTPUT_FIFO_19_DMWIDTH-1:0] m_axis_fifo_19_tdata,
    input m_axis_fifo_19_tready,
    output ap_fifo_oarg_19_full_n,
    input [C_OUTPUT_FIFO_19_WIDTH-1:0] ap_fifo_oarg_19_din,
    input ap_fifo_oarg_19_write,
    //output FIFO to AXI-Stream interface 20
    output m_axis_fifo_20_tlast,
    output m_axis_fifo_20_tvalid,
    output [C_OUTPUT_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tkeep,
    output [C_OUTPUT_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tstrb,
    output [C_OUTPUT_FIFO_20_DMWIDTH-1:0] m_axis_fifo_20_tdata,
    input m_axis_fifo_20_tready,
    output ap_fifo_oarg_20_full_n,
    input [C_OUTPUT_FIFO_20_WIDTH-1:0] ap_fifo_oarg_20_din,
    input ap_fifo_oarg_20_write,
    //output FIFO to AXI-Stream interface 21
    output m_axis_fifo_21_tlast,
    output m_axis_fifo_21_tvalid,
    output [C_OUTPUT_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tkeep,
    output [C_OUTPUT_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tstrb,
    output [C_OUTPUT_FIFO_21_DMWIDTH-1:0] m_axis_fifo_21_tdata,
    input m_axis_fifo_21_tready,
    output ap_fifo_oarg_21_full_n,
    input [C_OUTPUT_FIFO_21_WIDTH-1:0] ap_fifo_oarg_21_din,
    input ap_fifo_oarg_21_write,
    //output FIFO to AXI-Stream interface 22
    output m_axis_fifo_22_tlast,
    output m_axis_fifo_22_tvalid,
    output [C_OUTPUT_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tkeep,
    output [C_OUTPUT_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tstrb,
    output [C_OUTPUT_FIFO_22_DMWIDTH-1:0] m_axis_fifo_22_tdata,
    input m_axis_fifo_22_tready,
    output ap_fifo_oarg_22_full_n,
    input [C_OUTPUT_FIFO_22_WIDTH-1:0] ap_fifo_oarg_22_din,
    input ap_fifo_oarg_22_write,
    //output FIFO to AXI-Stream interface 23
    output m_axis_fifo_23_tlast,
    output m_axis_fifo_23_tvalid,
    output [C_OUTPUT_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tkeep,
    output [C_OUTPUT_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tstrb,
    output [C_OUTPUT_FIFO_23_DMWIDTH-1:0] m_axis_fifo_23_tdata,
    input m_axis_fifo_23_tready,
    output ap_fifo_oarg_23_full_n,
    input [C_OUTPUT_FIFO_23_WIDTH-1:0] ap_fifo_oarg_23_din,
    input ap_fifo_oarg_23_write,
    //output FIFO to AXI-Stream interface 24
    output m_axis_fifo_24_tlast,
    output m_axis_fifo_24_tvalid,
    output [C_OUTPUT_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tkeep,
    output [C_OUTPUT_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tstrb,
    output [C_OUTPUT_FIFO_24_DMWIDTH-1:0] m_axis_fifo_24_tdata,
    input m_axis_fifo_24_tready,
    output ap_fifo_oarg_24_full_n,
    input [C_OUTPUT_FIFO_24_WIDTH-1:0] ap_fifo_oarg_24_din,
    input ap_fifo_oarg_24_write,
    //output FIFO to AXI-Stream interface 25
    output m_axis_fifo_25_tlast,
    output m_axis_fifo_25_tvalid,
    output [C_OUTPUT_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tkeep,
    output [C_OUTPUT_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tstrb,
    output [C_OUTPUT_FIFO_25_DMWIDTH-1:0] m_axis_fifo_25_tdata,
    input m_axis_fifo_25_tready,
    output ap_fifo_oarg_25_full_n,
    input [C_OUTPUT_FIFO_25_WIDTH-1:0] ap_fifo_oarg_25_din,
    input ap_fifo_oarg_25_write,
    //output FIFO to AXI-Stream interface 26
    output m_axis_fifo_26_tlast,
    output m_axis_fifo_26_tvalid,
    output [C_OUTPUT_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tkeep,
    output [C_OUTPUT_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tstrb,
    output [C_OUTPUT_FIFO_26_DMWIDTH-1:0] m_axis_fifo_26_tdata,
    input m_axis_fifo_26_tready,
    output ap_fifo_oarg_26_full_n,
    input [C_OUTPUT_FIFO_26_WIDTH-1:0] ap_fifo_oarg_26_din,
    input ap_fifo_oarg_26_write,
    //output FIFO to AXI-Stream interface 27
    output m_axis_fifo_27_tlast,
    output m_axis_fifo_27_tvalid,
    output [C_OUTPUT_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tkeep,
    output [C_OUTPUT_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tstrb,
    output [C_OUTPUT_FIFO_27_DMWIDTH-1:0] m_axis_fifo_27_tdata,
    input m_axis_fifo_27_tready,
    output ap_fifo_oarg_27_full_n,
    input [C_OUTPUT_FIFO_27_WIDTH-1:0] ap_fifo_oarg_27_din,
    input ap_fifo_oarg_27_write,
    //output FIFO to AXI-Stream interface 28
    output m_axis_fifo_28_tlast,
    output m_axis_fifo_28_tvalid,
    output [C_OUTPUT_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tkeep,
    output [C_OUTPUT_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tstrb,
    output [C_OUTPUT_FIFO_28_DMWIDTH-1:0] m_axis_fifo_28_tdata,
    input m_axis_fifo_28_tready,
    output ap_fifo_oarg_28_full_n,
    input [C_OUTPUT_FIFO_28_WIDTH-1:0] ap_fifo_oarg_28_din,
    input ap_fifo_oarg_28_write,
    //output FIFO to AXI-Stream interface 29
    output m_axis_fifo_29_tlast,
    output m_axis_fifo_29_tvalid,
    output [C_OUTPUT_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tkeep,
    output [C_OUTPUT_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tstrb,
    output [C_OUTPUT_FIFO_29_DMWIDTH-1:0] m_axis_fifo_29_tdata,
    input m_axis_fifo_29_tready,
    output ap_fifo_oarg_29_full_n,
    input [C_OUTPUT_FIFO_29_WIDTH-1:0] ap_fifo_oarg_29_din,
    input ap_fifo_oarg_29_write,
    //output FIFO to AXI-Stream interface 30
    output m_axis_fifo_30_tlast,
    output m_axis_fifo_30_tvalid,
    output [C_OUTPUT_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tkeep,
    output [C_OUTPUT_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tstrb,
    output [C_OUTPUT_FIFO_30_DMWIDTH-1:0] m_axis_fifo_30_tdata,
    input m_axis_fifo_30_tready,
    output ap_fifo_oarg_30_full_n,
    input [C_OUTPUT_FIFO_30_WIDTH-1:0] ap_fifo_oarg_30_din,
    input ap_fifo_oarg_30_write,
    //output FIFO to AXI-Stream interface 31
    output m_axis_fifo_31_tlast,
    output m_axis_fifo_31_tvalid,
    output [C_OUTPUT_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tkeep,
    output [C_OUTPUT_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tstrb,
    output [C_OUTPUT_FIFO_31_DMWIDTH-1:0] m_axis_fifo_31_tdata,
    input m_axis_fifo_31_tready,
    output ap_fifo_oarg_31_full_n,
    input [C_OUTPUT_FIFO_31_WIDTH-1:0] ap_fifo_oarg_31_din,
    input ap_fifo_oarg_31_write,
    //output FIFO to AXI-Stream interface 32
    output m_axis_fifo_32_tlast,
    output m_axis_fifo_32_tvalid,
    output [C_OUTPUT_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tkeep,
    output [C_OUTPUT_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tstrb,
    output [C_OUTPUT_FIFO_32_DMWIDTH-1:0] m_axis_fifo_32_tdata,
    input m_axis_fifo_32_tready,
    output ap_fifo_oarg_32_full_n,
    input [C_OUTPUT_FIFO_32_WIDTH-1:0] ap_fifo_oarg_32_din,
    input ap_fifo_oarg_32_write,
    //output FIFO to AXI-Stream interface 33
    output m_axis_fifo_33_tlast,
    output m_axis_fifo_33_tvalid,
    output [C_OUTPUT_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tkeep,
    output [C_OUTPUT_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tstrb,
    output [C_OUTPUT_FIFO_33_DMWIDTH-1:0] m_axis_fifo_33_tdata,
    input m_axis_fifo_33_tready,
    output ap_fifo_oarg_33_full_n,
    input [C_OUTPUT_FIFO_33_WIDTH-1:0] ap_fifo_oarg_33_din,
    input ap_fifo_oarg_33_write,
    //output FIFO to AXI-Stream interface 34
    output m_axis_fifo_34_tlast,
    output m_axis_fifo_34_tvalid,
    output [C_OUTPUT_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tkeep,
    output [C_OUTPUT_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tstrb,
    output [C_OUTPUT_FIFO_34_DMWIDTH-1:0] m_axis_fifo_34_tdata,
    input m_axis_fifo_34_tready,
    output ap_fifo_oarg_34_full_n,
    input [C_OUTPUT_FIFO_34_WIDTH-1:0] ap_fifo_oarg_34_din,
    input ap_fifo_oarg_34_write,
    //output FIFO to AXI-Stream interface 35
    output m_axis_fifo_35_tlast,
    output m_axis_fifo_35_tvalid,
    output [C_OUTPUT_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tkeep,
    output [C_OUTPUT_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tstrb,
    output [C_OUTPUT_FIFO_35_DMWIDTH-1:0] m_axis_fifo_35_tdata,
    input m_axis_fifo_35_tready,
    output ap_fifo_oarg_35_full_n,
    input [C_OUTPUT_FIFO_35_WIDTH-1:0] ap_fifo_oarg_35_din,
    input ap_fifo_oarg_35_write,
    //output FIFO to AXI-Stream interface 36
    output m_axis_fifo_36_tlast,
    output m_axis_fifo_36_tvalid,
    output [C_OUTPUT_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tkeep,
    output [C_OUTPUT_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tstrb,
    output [C_OUTPUT_FIFO_36_DMWIDTH-1:0] m_axis_fifo_36_tdata,
    input m_axis_fifo_36_tready,
    output ap_fifo_oarg_36_full_n,
    input [C_OUTPUT_FIFO_36_WIDTH-1:0] ap_fifo_oarg_36_din,
    input ap_fifo_oarg_36_write,
    //output FIFO to AXI-Stream interface 37
    output m_axis_fifo_37_tlast,
    output m_axis_fifo_37_tvalid,
    output [C_OUTPUT_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tkeep,
    output [C_OUTPUT_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tstrb,
    output [C_OUTPUT_FIFO_37_DMWIDTH-1:0] m_axis_fifo_37_tdata,
    input m_axis_fifo_37_tready,
    output ap_fifo_oarg_37_full_n,
    input [C_OUTPUT_FIFO_37_WIDTH-1:0] ap_fifo_oarg_37_din,
    input ap_fifo_oarg_37_write,
    //output FIFO to AXI-Stream interface 38
    output m_axis_fifo_38_tlast,
    output m_axis_fifo_38_tvalid,
    output [C_OUTPUT_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tkeep,
    output [C_OUTPUT_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tstrb,
    output [C_OUTPUT_FIFO_38_DMWIDTH-1:0] m_axis_fifo_38_tdata,
    input m_axis_fifo_38_tready,
    output ap_fifo_oarg_38_full_n,
    input [C_OUTPUT_FIFO_38_WIDTH-1:0] ap_fifo_oarg_38_din,
    input ap_fifo_oarg_38_write,
    //output FIFO to AXI-Stream interface 39
    output m_axis_fifo_39_tlast,
    output m_axis_fifo_39_tvalid,
    output [C_OUTPUT_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tkeep,
    output [C_OUTPUT_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tstrb,
    output [C_OUTPUT_FIFO_39_DMWIDTH-1:0] m_axis_fifo_39_tdata,
    input m_axis_fifo_39_tready,
    output ap_fifo_oarg_39_full_n,
    input [C_OUTPUT_FIFO_39_WIDTH-1:0] ap_fifo_oarg_39_din,
    input ap_fifo_oarg_39_write,
    //output FIFO to AXI-Stream interface 40
    output m_axis_fifo_40_tlast,
    output m_axis_fifo_40_tvalid,
    output [C_OUTPUT_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tkeep,
    output [C_OUTPUT_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tstrb,
    output [C_OUTPUT_FIFO_40_DMWIDTH-1:0] m_axis_fifo_40_tdata,
    input m_axis_fifo_40_tready,
    output ap_fifo_oarg_40_full_n,
    input [C_OUTPUT_FIFO_40_WIDTH-1:0] ap_fifo_oarg_40_din,
    input ap_fifo_oarg_40_write,
    //output FIFO to AXI-Stream interface 41
    output m_axis_fifo_41_tlast,
    output m_axis_fifo_41_tvalid,
    output [C_OUTPUT_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tkeep,
    output [C_OUTPUT_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tstrb,
    output [C_OUTPUT_FIFO_41_DMWIDTH-1:0] m_axis_fifo_41_tdata,
    input m_axis_fifo_41_tready,
    output ap_fifo_oarg_41_full_n,
    input [C_OUTPUT_FIFO_41_WIDTH-1:0] ap_fifo_oarg_41_din,
    input ap_fifo_oarg_41_write,
    //output FIFO to AXI-Stream interface 42
    output m_axis_fifo_42_tlast,
    output m_axis_fifo_42_tvalid,
    output [C_OUTPUT_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tkeep,
    output [C_OUTPUT_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tstrb,
    output [C_OUTPUT_FIFO_42_DMWIDTH-1:0] m_axis_fifo_42_tdata,
    input m_axis_fifo_42_tready,
    output ap_fifo_oarg_42_full_n,
    input [C_OUTPUT_FIFO_42_WIDTH-1:0] ap_fifo_oarg_42_din,
    input ap_fifo_oarg_42_write,
    //output FIFO to AXI-Stream interface 43
    output m_axis_fifo_43_tlast,
    output m_axis_fifo_43_tvalid,
    output [C_OUTPUT_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tkeep,
    output [C_OUTPUT_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tstrb,
    output [C_OUTPUT_FIFO_43_DMWIDTH-1:0] m_axis_fifo_43_tdata,
    input m_axis_fifo_43_tready,
    output ap_fifo_oarg_43_full_n,
    input [C_OUTPUT_FIFO_43_WIDTH-1:0] ap_fifo_oarg_43_din,
    input ap_fifo_oarg_43_write,
    //output FIFO to AXI-Stream interface 44
    output m_axis_fifo_44_tlast,
    output m_axis_fifo_44_tvalid,
    output [C_OUTPUT_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tkeep,
    output [C_OUTPUT_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tstrb,
    output [C_OUTPUT_FIFO_44_DMWIDTH-1:0] m_axis_fifo_44_tdata,
    input m_axis_fifo_44_tready,
    output ap_fifo_oarg_44_full_n,
    input [C_OUTPUT_FIFO_44_WIDTH-1:0] ap_fifo_oarg_44_din,
    input ap_fifo_oarg_44_write,
    //output FIFO to AXI-Stream interface 45
    output m_axis_fifo_45_tlast,
    output m_axis_fifo_45_tvalid,
    output [C_OUTPUT_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tkeep,
    output [C_OUTPUT_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tstrb,
    output [C_OUTPUT_FIFO_45_DMWIDTH-1:0] m_axis_fifo_45_tdata,
    input m_axis_fifo_45_tready,
    output ap_fifo_oarg_45_full_n,
    input [C_OUTPUT_FIFO_45_WIDTH-1:0] ap_fifo_oarg_45_din,
    input ap_fifo_oarg_45_write,
    //output FIFO to AXI-Stream interface 46
    output m_axis_fifo_46_tlast,
    output m_axis_fifo_46_tvalid,
    output [C_OUTPUT_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tkeep,
    output [C_OUTPUT_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tstrb,
    output [C_OUTPUT_FIFO_46_DMWIDTH-1:0] m_axis_fifo_46_tdata,
    input m_axis_fifo_46_tready,
    output ap_fifo_oarg_46_full_n,
    input [C_OUTPUT_FIFO_46_WIDTH-1:0] ap_fifo_oarg_46_din,
    input ap_fifo_oarg_46_write,
    //output FIFO to AXI-Stream interface 47
    output m_axis_fifo_47_tlast,
    output m_axis_fifo_47_tvalid,
    output [C_OUTPUT_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tkeep,
    output [C_OUTPUT_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tstrb,
    output [C_OUTPUT_FIFO_47_DMWIDTH-1:0] m_axis_fifo_47_tdata,
    input m_axis_fifo_47_tready,
    output ap_fifo_oarg_47_full_n,
    input [C_OUTPUT_FIFO_47_WIDTH-1:0] ap_fifo_oarg_47_din,
    input ap_fifo_oarg_47_write,
    //output FIFO to AXI-Stream interface 48
    output m_axis_fifo_48_tlast,
    output m_axis_fifo_48_tvalid,
    output [C_OUTPUT_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tkeep,
    output [C_OUTPUT_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tstrb,
    output [C_OUTPUT_FIFO_48_DMWIDTH-1:0] m_axis_fifo_48_tdata,
    input m_axis_fifo_48_tready,
    output ap_fifo_oarg_48_full_n,
    input [C_OUTPUT_FIFO_48_WIDTH-1:0] ap_fifo_oarg_48_din,
    input ap_fifo_oarg_48_write,
    //output FIFO to AXI-Stream interface 49
    output m_axis_fifo_49_tlast,
    output m_axis_fifo_49_tvalid,
    output [C_OUTPUT_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tkeep,
    output [C_OUTPUT_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tstrb,
    output [C_OUTPUT_FIFO_49_DMWIDTH-1:0] m_axis_fifo_49_tdata,
    input m_axis_fifo_49_tready,
    output ap_fifo_oarg_49_full_n,
    input [C_OUTPUT_FIFO_49_WIDTH-1:0] ap_fifo_oarg_49_din,
    input ap_fifo_oarg_49_write,
    //output FIFO to AXI-Stream interface 50
    output m_axis_fifo_50_tlast,
    output m_axis_fifo_50_tvalid,
    output [C_OUTPUT_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tkeep,
    output [C_OUTPUT_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tstrb,
    output [C_OUTPUT_FIFO_50_DMWIDTH-1:0] m_axis_fifo_50_tdata,
    input m_axis_fifo_50_tready,
    output ap_fifo_oarg_50_full_n,
    input [C_OUTPUT_FIFO_50_WIDTH-1:0] ap_fifo_oarg_50_din,
    input ap_fifo_oarg_50_write,
    //output FIFO to AXI-Stream interface 51
    output m_axis_fifo_51_tlast,
    output m_axis_fifo_51_tvalid,
    output [C_OUTPUT_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tkeep,
    output [C_OUTPUT_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tstrb,
    output [C_OUTPUT_FIFO_51_DMWIDTH-1:0] m_axis_fifo_51_tdata,
    input m_axis_fifo_51_tready,
    output ap_fifo_oarg_51_full_n,
    input [C_OUTPUT_FIFO_51_WIDTH-1:0] ap_fifo_oarg_51_din,
    input ap_fifo_oarg_51_write,
    //output FIFO to AXI-Stream interface 52
    output m_axis_fifo_52_tlast,
    output m_axis_fifo_52_tvalid,
    output [C_OUTPUT_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tkeep,
    output [C_OUTPUT_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tstrb,
    output [C_OUTPUT_FIFO_52_DMWIDTH-1:0] m_axis_fifo_52_tdata,
    input m_axis_fifo_52_tready,
    output ap_fifo_oarg_52_full_n,
    input [C_OUTPUT_FIFO_52_WIDTH-1:0] ap_fifo_oarg_52_din,
    input ap_fifo_oarg_52_write,
    //output FIFO to AXI-Stream interface 53
    output m_axis_fifo_53_tlast,
    output m_axis_fifo_53_tvalid,
    output [C_OUTPUT_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tkeep,
    output [C_OUTPUT_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tstrb,
    output [C_OUTPUT_FIFO_53_DMWIDTH-1:0] m_axis_fifo_53_tdata,
    input m_axis_fifo_53_tready,
    output ap_fifo_oarg_53_full_n,
    input [C_OUTPUT_FIFO_53_WIDTH-1:0] ap_fifo_oarg_53_din,
    input ap_fifo_oarg_53_write,
    //output FIFO to AXI-Stream interface 54
    output m_axis_fifo_54_tlast,
    output m_axis_fifo_54_tvalid,
    output [C_OUTPUT_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tkeep,
    output [C_OUTPUT_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tstrb,
    output [C_OUTPUT_FIFO_54_DMWIDTH-1:0] m_axis_fifo_54_tdata,
    input m_axis_fifo_54_tready,
    output ap_fifo_oarg_54_full_n,
    input [C_OUTPUT_FIFO_54_WIDTH-1:0] ap_fifo_oarg_54_din,
    input ap_fifo_oarg_54_write,
    //output FIFO to AXI-Stream interface 55
    output m_axis_fifo_55_tlast,
    output m_axis_fifo_55_tvalid,
    output [C_OUTPUT_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tkeep,
    output [C_OUTPUT_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tstrb,
    output [C_OUTPUT_FIFO_55_DMWIDTH-1:0] m_axis_fifo_55_tdata,
    input m_axis_fifo_55_tready,
    output ap_fifo_oarg_55_full_n,
    input [C_OUTPUT_FIFO_55_WIDTH-1:0] ap_fifo_oarg_55_din,
    input ap_fifo_oarg_55_write,
    //output FIFO to AXI-Stream interface 56
    output m_axis_fifo_56_tlast,
    output m_axis_fifo_56_tvalid,
    output [C_OUTPUT_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tkeep,
    output [C_OUTPUT_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tstrb,
    output [C_OUTPUT_FIFO_56_DMWIDTH-1:0] m_axis_fifo_56_tdata,
    input m_axis_fifo_56_tready,
    output ap_fifo_oarg_56_full_n,
    input [C_OUTPUT_FIFO_56_WIDTH-1:0] ap_fifo_oarg_56_din,
    input ap_fifo_oarg_56_write,
    //output FIFO to AXI-Stream interface 57
    output m_axis_fifo_57_tlast,
    output m_axis_fifo_57_tvalid,
    output [C_OUTPUT_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tkeep,
    output [C_OUTPUT_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tstrb,
    output [C_OUTPUT_FIFO_57_DMWIDTH-1:0] m_axis_fifo_57_tdata,
    input m_axis_fifo_57_tready,
    output ap_fifo_oarg_57_full_n,
    input [C_OUTPUT_FIFO_57_WIDTH-1:0] ap_fifo_oarg_57_din,
    input ap_fifo_oarg_57_write,
    //output FIFO to AXI-Stream interface 58
    output m_axis_fifo_58_tlast,
    output m_axis_fifo_58_tvalid,
    output [C_OUTPUT_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tkeep,
    output [C_OUTPUT_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tstrb,
    output [C_OUTPUT_FIFO_58_DMWIDTH-1:0] m_axis_fifo_58_tdata,
    input m_axis_fifo_58_tready,
    output ap_fifo_oarg_58_full_n,
    input [C_OUTPUT_FIFO_58_WIDTH-1:0] ap_fifo_oarg_58_din,
    input ap_fifo_oarg_58_write,
    //output FIFO to AXI-Stream interface 59
    output m_axis_fifo_59_tlast,
    output m_axis_fifo_59_tvalid,
    output [C_OUTPUT_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tkeep,
    output [C_OUTPUT_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tstrb,
    output [C_OUTPUT_FIFO_59_DMWIDTH-1:0] m_axis_fifo_59_tdata,
    input m_axis_fifo_59_tready,
    output ap_fifo_oarg_59_full_n,
    input [C_OUTPUT_FIFO_59_WIDTH-1:0] ap_fifo_oarg_59_din,
    input ap_fifo_oarg_59_write,
    //output FIFO to AXI-Stream interface 60
    output m_axis_fifo_60_tlast,
    output m_axis_fifo_60_tvalid,
    output [C_OUTPUT_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tkeep,
    output [C_OUTPUT_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tstrb,
    output [C_OUTPUT_FIFO_60_DMWIDTH-1:0] m_axis_fifo_60_tdata,
    input m_axis_fifo_60_tready,
    output ap_fifo_oarg_60_full_n,
    input [C_OUTPUT_FIFO_60_WIDTH-1:0] ap_fifo_oarg_60_din,
    input ap_fifo_oarg_60_write,
    //output FIFO to AXI-Stream interface 61
    output m_axis_fifo_61_tlast,
    output m_axis_fifo_61_tvalid,
    output [C_OUTPUT_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tkeep,
    output [C_OUTPUT_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tstrb,
    output [C_OUTPUT_FIFO_61_DMWIDTH-1:0] m_axis_fifo_61_tdata,
    input m_axis_fifo_61_tready,
    output ap_fifo_oarg_61_full_n,
    input [C_OUTPUT_FIFO_61_WIDTH-1:0] ap_fifo_oarg_61_din,
    input ap_fifo_oarg_61_write,
    //output FIFO to AXI-Stream interface 62
    output m_axis_fifo_62_tlast,
    output m_axis_fifo_62_tvalid,
    output [C_OUTPUT_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tkeep,
    output [C_OUTPUT_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tstrb,
    output [C_OUTPUT_FIFO_62_DMWIDTH-1:0] m_axis_fifo_62_tdata,
    input m_axis_fifo_62_tready,
    output ap_fifo_oarg_62_full_n,
    input [C_OUTPUT_FIFO_62_WIDTH-1:0] ap_fifo_oarg_62_din,
    input ap_fifo_oarg_62_write,
    //output FIFO to AXI-Stream interface 63
    output m_axis_fifo_63_tlast,
    output m_axis_fifo_63_tvalid,
    output [C_OUTPUT_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tkeep,
    output [C_OUTPUT_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tstrb,
    output [C_OUTPUT_FIFO_63_DMWIDTH-1:0] m_axis_fifo_63_tdata,
    input m_axis_fifo_63_tready,
    output ap_fifo_oarg_63_full_n,
    input [C_OUTPUT_FIFO_63_WIDTH-1:0] ap_fifo_oarg_63_din,
    input ap_fifo_oarg_63_write,
    //output FIFO to AXI-Stream interface 64
    output m_axis_fifo_64_tlast,
    output m_axis_fifo_64_tvalid,
    output [C_OUTPUT_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tkeep,
    output [C_OUTPUT_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tstrb,
    output [C_OUTPUT_FIFO_64_DMWIDTH-1:0] m_axis_fifo_64_tdata,
    input m_axis_fifo_64_tready,
    output ap_fifo_oarg_64_full_n,
    input [C_OUTPUT_FIFO_64_WIDTH-1:0] ap_fifo_oarg_64_din,
    input ap_fifo_oarg_64_write,
    //output FIFO to AXI-Stream interface 65
    output m_axis_fifo_65_tlast,
    output m_axis_fifo_65_tvalid,
    output [C_OUTPUT_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tkeep,
    output [C_OUTPUT_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tstrb,
    output [C_OUTPUT_FIFO_65_DMWIDTH-1:0] m_axis_fifo_65_tdata,
    input m_axis_fifo_65_tready,
    output ap_fifo_oarg_65_full_n,
    input [C_OUTPUT_FIFO_65_WIDTH-1:0] ap_fifo_oarg_65_din,
    input ap_fifo_oarg_65_write,
    //output FIFO to AXI-Stream interface 66
    output m_axis_fifo_66_tlast,
    output m_axis_fifo_66_tvalid,
    output [C_OUTPUT_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tkeep,
    output [C_OUTPUT_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tstrb,
    output [C_OUTPUT_FIFO_66_DMWIDTH-1:0] m_axis_fifo_66_tdata,
    input m_axis_fifo_66_tready,
    output ap_fifo_oarg_66_full_n,
    input [C_OUTPUT_FIFO_66_WIDTH-1:0] ap_fifo_oarg_66_din,
    input ap_fifo_oarg_66_write,
    //output FIFO to AXI-Stream interface 67
    output m_axis_fifo_67_tlast,
    output m_axis_fifo_67_tvalid,
    output [C_OUTPUT_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tkeep,
    output [C_OUTPUT_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tstrb,
    output [C_OUTPUT_FIFO_67_DMWIDTH-1:0] m_axis_fifo_67_tdata,
    input m_axis_fifo_67_tready,
    output ap_fifo_oarg_67_full_n,
    input [C_OUTPUT_FIFO_67_WIDTH-1:0] ap_fifo_oarg_67_din,
    input ap_fifo_oarg_67_write,
    //output FIFO to AXI-Stream interface 68
    output m_axis_fifo_68_tlast,
    output m_axis_fifo_68_tvalid,
    output [C_OUTPUT_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tkeep,
    output [C_OUTPUT_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tstrb,
    output [C_OUTPUT_FIFO_68_DMWIDTH-1:0] m_axis_fifo_68_tdata,
    input m_axis_fifo_68_tready,
    output ap_fifo_oarg_68_full_n,
    input [C_OUTPUT_FIFO_68_WIDTH-1:0] ap_fifo_oarg_68_din,
    input ap_fifo_oarg_68_write,
    //output FIFO to AXI-Stream interface 69
    output m_axis_fifo_69_tlast,
    output m_axis_fifo_69_tvalid,
    output [C_OUTPUT_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tkeep,
    output [C_OUTPUT_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tstrb,
    output [C_OUTPUT_FIFO_69_DMWIDTH-1:0] m_axis_fifo_69_tdata,
    input m_axis_fifo_69_tready,
    output ap_fifo_oarg_69_full_n,
    input [C_OUTPUT_FIFO_69_WIDTH-1:0] ap_fifo_oarg_69_din,
    input ap_fifo_oarg_69_write,
    //output FIFO to AXI-Stream interface 70
    output m_axis_fifo_70_tlast,
    output m_axis_fifo_70_tvalid,
    output [C_OUTPUT_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tkeep,
    output [C_OUTPUT_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tstrb,
    output [C_OUTPUT_FIFO_70_DMWIDTH-1:0] m_axis_fifo_70_tdata,
    input m_axis_fifo_70_tready,
    output ap_fifo_oarg_70_full_n,
    input [C_OUTPUT_FIFO_70_WIDTH-1:0] ap_fifo_oarg_70_din,
    input ap_fifo_oarg_70_write,
    //output FIFO to AXI-Stream interface 71
    output m_axis_fifo_71_tlast,
    output m_axis_fifo_71_tvalid,
    output [C_OUTPUT_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tkeep,
    output [C_OUTPUT_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tstrb,
    output [C_OUTPUT_FIFO_71_DMWIDTH-1:0] m_axis_fifo_71_tdata,
    input m_axis_fifo_71_tready,
    output ap_fifo_oarg_71_full_n,
    input [C_OUTPUT_FIFO_71_WIDTH-1:0] ap_fifo_oarg_71_din,
    input ap_fifo_oarg_71_write,
    //output FIFO to AXI-Stream interface 72
    output m_axis_fifo_72_tlast,
    output m_axis_fifo_72_tvalid,
    output [C_OUTPUT_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tkeep,
    output [C_OUTPUT_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tstrb,
    output [C_OUTPUT_FIFO_72_DMWIDTH-1:0] m_axis_fifo_72_tdata,
    input m_axis_fifo_72_tready,
    output ap_fifo_oarg_72_full_n,
    input [C_OUTPUT_FIFO_72_WIDTH-1:0] ap_fifo_oarg_72_din,
    input ap_fifo_oarg_72_write,
    //output FIFO to AXI-Stream interface 73
    output m_axis_fifo_73_tlast,
    output m_axis_fifo_73_tvalid,
    output [C_OUTPUT_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tkeep,
    output [C_OUTPUT_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tstrb,
    output [C_OUTPUT_FIFO_73_DMWIDTH-1:0] m_axis_fifo_73_tdata,
    input m_axis_fifo_73_tready,
    output ap_fifo_oarg_73_full_n,
    input [C_OUTPUT_FIFO_73_WIDTH-1:0] ap_fifo_oarg_73_din,
    input ap_fifo_oarg_73_write,
    //output FIFO to AXI-Stream interface 74
    output m_axis_fifo_74_tlast,
    output m_axis_fifo_74_tvalid,
    output [C_OUTPUT_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tkeep,
    output [C_OUTPUT_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tstrb,
    output [C_OUTPUT_FIFO_74_DMWIDTH-1:0] m_axis_fifo_74_tdata,
    input m_axis_fifo_74_tready,
    output ap_fifo_oarg_74_full_n,
    input [C_OUTPUT_FIFO_74_WIDTH-1:0] ap_fifo_oarg_74_din,
    input ap_fifo_oarg_74_write,
    //output FIFO to AXI-Stream interface 75
    output m_axis_fifo_75_tlast,
    output m_axis_fifo_75_tvalid,
    output [C_OUTPUT_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tkeep,
    output [C_OUTPUT_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tstrb,
    output [C_OUTPUT_FIFO_75_DMWIDTH-1:0] m_axis_fifo_75_tdata,
    input m_axis_fifo_75_tready,
    output ap_fifo_oarg_75_full_n,
    input [C_OUTPUT_FIFO_75_WIDTH-1:0] ap_fifo_oarg_75_din,
    input ap_fifo_oarg_75_write,
    //output FIFO to AXI-Stream interface 76
    output m_axis_fifo_76_tlast,
    output m_axis_fifo_76_tvalid,
    output [C_OUTPUT_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tkeep,
    output [C_OUTPUT_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tstrb,
    output [C_OUTPUT_FIFO_76_DMWIDTH-1:0] m_axis_fifo_76_tdata,
    input m_axis_fifo_76_tready,
    output ap_fifo_oarg_76_full_n,
    input [C_OUTPUT_FIFO_76_WIDTH-1:0] ap_fifo_oarg_76_din,
    input ap_fifo_oarg_76_write,
    //output FIFO to AXI-Stream interface 77
    output m_axis_fifo_77_tlast,
    output m_axis_fifo_77_tvalid,
    output [C_OUTPUT_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tkeep,
    output [C_OUTPUT_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tstrb,
    output [C_OUTPUT_FIFO_77_DMWIDTH-1:0] m_axis_fifo_77_tdata,
    input m_axis_fifo_77_tready,
    output ap_fifo_oarg_77_full_n,
    input [C_OUTPUT_FIFO_77_WIDTH-1:0] ap_fifo_oarg_77_din,
    input ap_fifo_oarg_77_write,
    //output FIFO to AXI-Stream interface 78
    output m_axis_fifo_78_tlast,
    output m_axis_fifo_78_tvalid,
    output [C_OUTPUT_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tkeep,
    output [C_OUTPUT_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tstrb,
    output [C_OUTPUT_FIFO_78_DMWIDTH-1:0] m_axis_fifo_78_tdata,
    input m_axis_fifo_78_tready,
    output ap_fifo_oarg_78_full_n,
    input [C_OUTPUT_FIFO_78_WIDTH-1:0] ap_fifo_oarg_78_din,
    input ap_fifo_oarg_78_write,
    //output FIFO to AXI-Stream interface 79
    output m_axis_fifo_79_tlast,
    output m_axis_fifo_79_tvalid,
    output [C_OUTPUT_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tkeep,
    output [C_OUTPUT_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tstrb,
    output [C_OUTPUT_FIFO_79_DMWIDTH-1:0] m_axis_fifo_79_tdata,
    input m_axis_fifo_79_tready,
    output ap_fifo_oarg_79_full_n,
    input [C_OUTPUT_FIFO_79_WIDTH-1:0] ap_fifo_oarg_79_din,
    input ap_fifo_oarg_79_write,
    //output FIFO to AXI-Stream interface 80
    output m_axis_fifo_80_tlast,
    output m_axis_fifo_80_tvalid,
    output [C_OUTPUT_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tkeep,
    output [C_OUTPUT_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tstrb,
    output [C_OUTPUT_FIFO_80_DMWIDTH-1:0] m_axis_fifo_80_tdata,
    input m_axis_fifo_80_tready,
    output ap_fifo_oarg_80_full_n,
    input [C_OUTPUT_FIFO_80_WIDTH-1:0] ap_fifo_oarg_80_din,
    input ap_fifo_oarg_80_write,
    //output FIFO to AXI-Stream interface 81
    output m_axis_fifo_81_tlast,
    output m_axis_fifo_81_tvalid,
    output [C_OUTPUT_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tkeep,
    output [C_OUTPUT_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tstrb,
    output [C_OUTPUT_FIFO_81_DMWIDTH-1:0] m_axis_fifo_81_tdata,
    input m_axis_fifo_81_tready,
    output ap_fifo_oarg_81_full_n,
    input [C_OUTPUT_FIFO_81_WIDTH-1:0] ap_fifo_oarg_81_din,
    input ap_fifo_oarg_81_write,
    //output FIFO to AXI-Stream interface 82
    output m_axis_fifo_82_tlast,
    output m_axis_fifo_82_tvalid,
    output [C_OUTPUT_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tkeep,
    output [C_OUTPUT_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tstrb,
    output [C_OUTPUT_FIFO_82_DMWIDTH-1:0] m_axis_fifo_82_tdata,
    input m_axis_fifo_82_tready,
    output ap_fifo_oarg_82_full_n,
    input [C_OUTPUT_FIFO_82_WIDTH-1:0] ap_fifo_oarg_82_din,
    input ap_fifo_oarg_82_write,
    //output FIFO to AXI-Stream interface 83
    output m_axis_fifo_83_tlast,
    output m_axis_fifo_83_tvalid,
    output [C_OUTPUT_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tkeep,
    output [C_OUTPUT_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tstrb,
    output [C_OUTPUT_FIFO_83_DMWIDTH-1:0] m_axis_fifo_83_tdata,
    input m_axis_fifo_83_tready,
    output ap_fifo_oarg_83_full_n,
    input [C_OUTPUT_FIFO_83_WIDTH-1:0] ap_fifo_oarg_83_din,
    input ap_fifo_oarg_83_write,
    //output FIFO to AXI-Stream interface 84
    output m_axis_fifo_84_tlast,
    output m_axis_fifo_84_tvalid,
    output [C_OUTPUT_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tkeep,
    output [C_OUTPUT_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tstrb,
    output [C_OUTPUT_FIFO_84_DMWIDTH-1:0] m_axis_fifo_84_tdata,
    input m_axis_fifo_84_tready,
    output ap_fifo_oarg_84_full_n,
    input [C_OUTPUT_FIFO_84_WIDTH-1:0] ap_fifo_oarg_84_din,
    input ap_fifo_oarg_84_write,
    //output FIFO to AXI-Stream interface 85
    output m_axis_fifo_85_tlast,
    output m_axis_fifo_85_tvalid,
    output [C_OUTPUT_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tkeep,
    output [C_OUTPUT_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tstrb,
    output [C_OUTPUT_FIFO_85_DMWIDTH-1:0] m_axis_fifo_85_tdata,
    input m_axis_fifo_85_tready,
    output ap_fifo_oarg_85_full_n,
    input [C_OUTPUT_FIFO_85_WIDTH-1:0] ap_fifo_oarg_85_din,
    input ap_fifo_oarg_85_write,
    //output FIFO to AXI-Stream interface 86
    output m_axis_fifo_86_tlast,
    output m_axis_fifo_86_tvalid,
    output [C_OUTPUT_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tkeep,
    output [C_OUTPUT_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tstrb,
    output [C_OUTPUT_FIFO_86_DMWIDTH-1:0] m_axis_fifo_86_tdata,
    input m_axis_fifo_86_tready,
    output ap_fifo_oarg_86_full_n,
    input [C_OUTPUT_FIFO_86_WIDTH-1:0] ap_fifo_oarg_86_din,
    input ap_fifo_oarg_86_write,
    //output FIFO to AXI-Stream interface 87
    output m_axis_fifo_87_tlast,
    output m_axis_fifo_87_tvalid,
    output [C_OUTPUT_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tkeep,
    output [C_OUTPUT_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tstrb,
    output [C_OUTPUT_FIFO_87_DMWIDTH-1:0] m_axis_fifo_87_tdata,
    input m_axis_fifo_87_tready,
    output ap_fifo_oarg_87_full_n,
    input [C_OUTPUT_FIFO_87_WIDTH-1:0] ap_fifo_oarg_87_din,
    input ap_fifo_oarg_87_write,
    //output FIFO to AXI-Stream interface 88
    output m_axis_fifo_88_tlast,
    output m_axis_fifo_88_tvalid,
    output [C_OUTPUT_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tkeep,
    output [C_OUTPUT_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tstrb,
    output [C_OUTPUT_FIFO_88_DMWIDTH-1:0] m_axis_fifo_88_tdata,
    input m_axis_fifo_88_tready,
    output ap_fifo_oarg_88_full_n,
    input [C_OUTPUT_FIFO_88_WIDTH-1:0] ap_fifo_oarg_88_din,
    input ap_fifo_oarg_88_write,
    //output FIFO to AXI-Stream interface 89
    output m_axis_fifo_89_tlast,
    output m_axis_fifo_89_tvalid,
    output [C_OUTPUT_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tkeep,
    output [C_OUTPUT_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tstrb,
    output [C_OUTPUT_FIFO_89_DMWIDTH-1:0] m_axis_fifo_89_tdata,
    input m_axis_fifo_89_tready,
    output ap_fifo_oarg_89_full_n,
    input [C_OUTPUT_FIFO_89_WIDTH-1:0] ap_fifo_oarg_89_din,
    input ap_fifo_oarg_89_write,
    //output FIFO to AXI-Stream interface 90
    output m_axis_fifo_90_tlast,
    output m_axis_fifo_90_tvalid,
    output [C_OUTPUT_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tkeep,
    output [C_OUTPUT_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tstrb,
    output [C_OUTPUT_FIFO_90_DMWIDTH-1:0] m_axis_fifo_90_tdata,
    input m_axis_fifo_90_tready,
    output ap_fifo_oarg_90_full_n,
    input [C_OUTPUT_FIFO_90_WIDTH-1:0] ap_fifo_oarg_90_din,
    input ap_fifo_oarg_90_write,
    //output FIFO to AXI-Stream interface 91
    output m_axis_fifo_91_tlast,
    output m_axis_fifo_91_tvalid,
    output [C_OUTPUT_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tkeep,
    output [C_OUTPUT_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tstrb,
    output [C_OUTPUT_FIFO_91_DMWIDTH-1:0] m_axis_fifo_91_tdata,
    input m_axis_fifo_91_tready,
    output ap_fifo_oarg_91_full_n,
    input [C_OUTPUT_FIFO_91_WIDTH-1:0] ap_fifo_oarg_91_din,
    input ap_fifo_oarg_91_write,
    //output FIFO to AXI-Stream interface 92
    output m_axis_fifo_92_tlast,
    output m_axis_fifo_92_tvalid,
    output [C_OUTPUT_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tkeep,
    output [C_OUTPUT_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tstrb,
    output [C_OUTPUT_FIFO_92_DMWIDTH-1:0] m_axis_fifo_92_tdata,
    input m_axis_fifo_92_tready,
    output ap_fifo_oarg_92_full_n,
    input [C_OUTPUT_FIFO_92_WIDTH-1:0] ap_fifo_oarg_92_din,
    input ap_fifo_oarg_92_write,
    //output FIFO to AXI-Stream interface 93
    output m_axis_fifo_93_tlast,
    output m_axis_fifo_93_tvalid,
    output [C_OUTPUT_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tkeep,
    output [C_OUTPUT_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tstrb,
    output [C_OUTPUT_FIFO_93_DMWIDTH-1:0] m_axis_fifo_93_tdata,
    input m_axis_fifo_93_tready,
    output ap_fifo_oarg_93_full_n,
    input [C_OUTPUT_FIFO_93_WIDTH-1:0] ap_fifo_oarg_93_din,
    input ap_fifo_oarg_93_write,
    //output FIFO to AXI-Stream interface 94
    output m_axis_fifo_94_tlast,
    output m_axis_fifo_94_tvalid,
    output [C_OUTPUT_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tkeep,
    output [C_OUTPUT_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tstrb,
    output [C_OUTPUT_FIFO_94_DMWIDTH-1:0] m_axis_fifo_94_tdata,
    input m_axis_fifo_94_tready,
    output ap_fifo_oarg_94_full_n,
    input [C_OUTPUT_FIFO_94_WIDTH-1:0] ap_fifo_oarg_94_din,
    input ap_fifo_oarg_94_write,
    //output FIFO to AXI-Stream interface 95
    output m_axis_fifo_95_tlast,
    output m_axis_fifo_95_tvalid,
    output [C_OUTPUT_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tkeep,
    output [C_OUTPUT_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tstrb,
    output [C_OUTPUT_FIFO_95_DMWIDTH-1:0] m_axis_fifo_95_tdata,
    input m_axis_fifo_95_tready,
    output ap_fifo_oarg_95_full_n,
    input [C_OUTPUT_FIFO_95_WIDTH-1:0] ap_fifo_oarg_95_din,
    input ap_fifo_oarg_95_write,
    //output FIFO to AXI-Stream interface 96
    output m_axis_fifo_96_tlast,
    output m_axis_fifo_96_tvalid,
    output [C_OUTPUT_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tkeep,
    output [C_OUTPUT_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tstrb,
    output [C_OUTPUT_FIFO_96_DMWIDTH-1:0] m_axis_fifo_96_tdata,
    input m_axis_fifo_96_tready,
    output ap_fifo_oarg_96_full_n,
    input [C_OUTPUT_FIFO_96_WIDTH-1:0] ap_fifo_oarg_96_din,
    input ap_fifo_oarg_96_write,
    //output FIFO to AXI-Stream interface 97
    output m_axis_fifo_97_tlast,
    output m_axis_fifo_97_tvalid,
    output [C_OUTPUT_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tkeep,
    output [C_OUTPUT_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tstrb,
    output [C_OUTPUT_FIFO_97_DMWIDTH-1:0] m_axis_fifo_97_tdata,
    input m_axis_fifo_97_tready,
    output ap_fifo_oarg_97_full_n,
    input [C_OUTPUT_FIFO_97_WIDTH-1:0] ap_fifo_oarg_97_din,
    input ap_fifo_oarg_97_write,
    //output FIFO to AXI-Stream interface 98
    output m_axis_fifo_98_tlast,
    output m_axis_fifo_98_tvalid,
    output [C_OUTPUT_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tkeep,
    output [C_OUTPUT_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tstrb,
    output [C_OUTPUT_FIFO_98_DMWIDTH-1:0] m_axis_fifo_98_tdata,
    input m_axis_fifo_98_tready,
    output ap_fifo_oarg_98_full_n,
    input [C_OUTPUT_FIFO_98_WIDTH-1:0] ap_fifo_oarg_98_din,
    input ap_fifo_oarg_98_write,
    //output FIFO to AXI-Stream interface 99
    output m_axis_fifo_99_tlast,
    output m_axis_fifo_99_tvalid,
    output [C_OUTPUT_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tkeep,
    output [C_OUTPUT_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tstrb,
    output [C_OUTPUT_FIFO_99_DMWIDTH-1:0] m_axis_fifo_99_tdata,
    input m_axis_fifo_99_tready,
    output ap_fifo_oarg_99_full_n,
    input [C_OUTPUT_FIFO_99_WIDTH-1:0] ap_fifo_oarg_99_din,
    input ap_fifo_oarg_99_write,
    //output FIFO to AXI-Stream interface 100
    output m_axis_fifo_100_tlast,
    output m_axis_fifo_100_tvalid,
    output [C_OUTPUT_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tkeep,
    output [C_OUTPUT_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tstrb,
    output [C_OUTPUT_FIFO_100_DMWIDTH-1:0] m_axis_fifo_100_tdata,
    input m_axis_fifo_100_tready,
    output ap_fifo_oarg_100_full_n,
    input [C_OUTPUT_FIFO_100_WIDTH-1:0] ap_fifo_oarg_100_din,
    input ap_fifo_oarg_100_write,
    //output FIFO to AXI-Stream interface 101
    output m_axis_fifo_101_tlast,
    output m_axis_fifo_101_tvalid,
    output [C_OUTPUT_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tkeep,
    output [C_OUTPUT_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tstrb,
    output [C_OUTPUT_FIFO_101_DMWIDTH-1:0] m_axis_fifo_101_tdata,
    input m_axis_fifo_101_tready,
    output ap_fifo_oarg_101_full_n,
    input [C_OUTPUT_FIFO_101_WIDTH-1:0] ap_fifo_oarg_101_din,
    input ap_fifo_oarg_101_write,
    //output FIFO to AXI-Stream interface 102
    output m_axis_fifo_102_tlast,
    output m_axis_fifo_102_tvalid,
    output [C_OUTPUT_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tkeep,
    output [C_OUTPUT_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tstrb,
    output [C_OUTPUT_FIFO_102_DMWIDTH-1:0] m_axis_fifo_102_tdata,
    input m_axis_fifo_102_tready,
    output ap_fifo_oarg_102_full_n,
    input [C_OUTPUT_FIFO_102_WIDTH-1:0] ap_fifo_oarg_102_din,
    input ap_fifo_oarg_102_write,
    //output FIFO to AXI-Stream interface 103
    output m_axis_fifo_103_tlast,
    output m_axis_fifo_103_tvalid,
    output [C_OUTPUT_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tkeep,
    output [C_OUTPUT_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tstrb,
    output [C_OUTPUT_FIFO_103_DMWIDTH-1:0] m_axis_fifo_103_tdata,
    input m_axis_fifo_103_tready,
    output ap_fifo_oarg_103_full_n,
    input [C_OUTPUT_FIFO_103_WIDTH-1:0] ap_fifo_oarg_103_din,
    input ap_fifo_oarg_103_write,
    //output FIFO to AXI-Stream interface 104
    output m_axis_fifo_104_tlast,
    output m_axis_fifo_104_tvalid,
    output [C_OUTPUT_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tkeep,
    output [C_OUTPUT_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tstrb,
    output [C_OUTPUT_FIFO_104_DMWIDTH-1:0] m_axis_fifo_104_tdata,
    input m_axis_fifo_104_tready,
    output ap_fifo_oarg_104_full_n,
    input [C_OUTPUT_FIFO_104_WIDTH-1:0] ap_fifo_oarg_104_din,
    input ap_fifo_oarg_104_write,
    //output FIFO to AXI-Stream interface 105
    output m_axis_fifo_105_tlast,
    output m_axis_fifo_105_tvalid,
    output [C_OUTPUT_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tkeep,
    output [C_OUTPUT_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tstrb,
    output [C_OUTPUT_FIFO_105_DMWIDTH-1:0] m_axis_fifo_105_tdata,
    input m_axis_fifo_105_tready,
    output ap_fifo_oarg_105_full_n,
    input [C_OUTPUT_FIFO_105_WIDTH-1:0] ap_fifo_oarg_105_din,
    input ap_fifo_oarg_105_write,
    //output FIFO to AXI-Stream interface 106
    output m_axis_fifo_106_tlast,
    output m_axis_fifo_106_tvalid,
    output [C_OUTPUT_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tkeep,
    output [C_OUTPUT_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tstrb,
    output [C_OUTPUT_FIFO_106_DMWIDTH-1:0] m_axis_fifo_106_tdata,
    input m_axis_fifo_106_tready,
    output ap_fifo_oarg_106_full_n,
    input [C_OUTPUT_FIFO_106_WIDTH-1:0] ap_fifo_oarg_106_din,
    input ap_fifo_oarg_106_write,
    //output FIFO to AXI-Stream interface 107
    output m_axis_fifo_107_tlast,
    output m_axis_fifo_107_tvalid,
    output [C_OUTPUT_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tkeep,
    output [C_OUTPUT_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tstrb,
    output [C_OUTPUT_FIFO_107_DMWIDTH-1:0] m_axis_fifo_107_tdata,
    input m_axis_fifo_107_tready,
    output ap_fifo_oarg_107_full_n,
    input [C_OUTPUT_FIFO_107_WIDTH-1:0] ap_fifo_oarg_107_din,
    input ap_fifo_oarg_107_write,
    //output FIFO to AXI-Stream interface 108
    output m_axis_fifo_108_tlast,
    output m_axis_fifo_108_tvalid,
    output [C_OUTPUT_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tkeep,
    output [C_OUTPUT_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tstrb,
    output [C_OUTPUT_FIFO_108_DMWIDTH-1:0] m_axis_fifo_108_tdata,
    input m_axis_fifo_108_tready,
    output ap_fifo_oarg_108_full_n,
    input [C_OUTPUT_FIFO_108_WIDTH-1:0] ap_fifo_oarg_108_din,
    input ap_fifo_oarg_108_write,
    //output FIFO to AXI-Stream interface 109
    output m_axis_fifo_109_tlast,
    output m_axis_fifo_109_tvalid,
    output [C_OUTPUT_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tkeep,
    output [C_OUTPUT_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tstrb,
    output [C_OUTPUT_FIFO_109_DMWIDTH-1:0] m_axis_fifo_109_tdata,
    input m_axis_fifo_109_tready,
    output ap_fifo_oarg_109_full_n,
    input [C_OUTPUT_FIFO_109_WIDTH-1:0] ap_fifo_oarg_109_din,
    input ap_fifo_oarg_109_write,
    //output FIFO to AXI-Stream interface 110
    output m_axis_fifo_110_tlast,
    output m_axis_fifo_110_tvalid,
    output [C_OUTPUT_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tkeep,
    output [C_OUTPUT_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tstrb,
    output [C_OUTPUT_FIFO_110_DMWIDTH-1:0] m_axis_fifo_110_tdata,
    input m_axis_fifo_110_tready,
    output ap_fifo_oarg_110_full_n,
    input [C_OUTPUT_FIFO_110_WIDTH-1:0] ap_fifo_oarg_110_din,
    input ap_fifo_oarg_110_write,
    //output FIFO to AXI-Stream interface 111
    output m_axis_fifo_111_tlast,
    output m_axis_fifo_111_tvalid,
    output [C_OUTPUT_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tkeep,
    output [C_OUTPUT_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tstrb,
    output [C_OUTPUT_FIFO_111_DMWIDTH-1:0] m_axis_fifo_111_tdata,
    input m_axis_fifo_111_tready,
    output ap_fifo_oarg_111_full_n,
    input [C_OUTPUT_FIFO_111_WIDTH-1:0] ap_fifo_oarg_111_din,
    input ap_fifo_oarg_111_write,
    //output FIFO to AXI-Stream interface 112
    output m_axis_fifo_112_tlast,
    output m_axis_fifo_112_tvalid,
    output [C_OUTPUT_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tkeep,
    output [C_OUTPUT_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tstrb,
    output [C_OUTPUT_FIFO_112_DMWIDTH-1:0] m_axis_fifo_112_tdata,
    input m_axis_fifo_112_tready,
    output ap_fifo_oarg_112_full_n,
    input [C_OUTPUT_FIFO_112_WIDTH-1:0] ap_fifo_oarg_112_din,
    input ap_fifo_oarg_112_write,
    //output FIFO to AXI-Stream interface 113
    output m_axis_fifo_113_tlast,
    output m_axis_fifo_113_tvalid,
    output [C_OUTPUT_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tkeep,
    output [C_OUTPUT_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tstrb,
    output [C_OUTPUT_FIFO_113_DMWIDTH-1:0] m_axis_fifo_113_tdata,
    input m_axis_fifo_113_tready,
    output ap_fifo_oarg_113_full_n,
    input [C_OUTPUT_FIFO_113_WIDTH-1:0] ap_fifo_oarg_113_din,
    input ap_fifo_oarg_113_write,
    //output FIFO to AXI-Stream interface 114
    output m_axis_fifo_114_tlast,
    output m_axis_fifo_114_tvalid,
    output [C_OUTPUT_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tkeep,
    output [C_OUTPUT_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tstrb,
    output [C_OUTPUT_FIFO_114_DMWIDTH-1:0] m_axis_fifo_114_tdata,
    input m_axis_fifo_114_tready,
    output ap_fifo_oarg_114_full_n,
    input [C_OUTPUT_FIFO_114_WIDTH-1:0] ap_fifo_oarg_114_din,
    input ap_fifo_oarg_114_write,
    //output FIFO to AXI-Stream interface 115
    output m_axis_fifo_115_tlast,
    output m_axis_fifo_115_tvalid,
    output [C_OUTPUT_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tkeep,
    output [C_OUTPUT_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tstrb,
    output [C_OUTPUT_FIFO_115_DMWIDTH-1:0] m_axis_fifo_115_tdata,
    input m_axis_fifo_115_tready,
    output ap_fifo_oarg_115_full_n,
    input [C_OUTPUT_FIFO_115_WIDTH-1:0] ap_fifo_oarg_115_din,
    input ap_fifo_oarg_115_write,
    //output FIFO to AXI-Stream interface 116
    output m_axis_fifo_116_tlast,
    output m_axis_fifo_116_tvalid,
    output [C_OUTPUT_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tkeep,
    output [C_OUTPUT_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tstrb,
    output [C_OUTPUT_FIFO_116_DMWIDTH-1:0] m_axis_fifo_116_tdata,
    input m_axis_fifo_116_tready,
    output ap_fifo_oarg_116_full_n,
    input [C_OUTPUT_FIFO_116_WIDTH-1:0] ap_fifo_oarg_116_din,
    input ap_fifo_oarg_116_write,
    //output FIFO to AXI-Stream interface 117
    output m_axis_fifo_117_tlast,
    output m_axis_fifo_117_tvalid,
    output [C_OUTPUT_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tkeep,
    output [C_OUTPUT_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tstrb,
    output [C_OUTPUT_FIFO_117_DMWIDTH-1:0] m_axis_fifo_117_tdata,
    input m_axis_fifo_117_tready,
    output ap_fifo_oarg_117_full_n,
    input [C_OUTPUT_FIFO_117_WIDTH-1:0] ap_fifo_oarg_117_din,
    input ap_fifo_oarg_117_write,
    //output FIFO to AXI-Stream interface 118
    output m_axis_fifo_118_tlast,
    output m_axis_fifo_118_tvalid,
    output [C_OUTPUT_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tkeep,
    output [C_OUTPUT_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tstrb,
    output [C_OUTPUT_FIFO_118_DMWIDTH-1:0] m_axis_fifo_118_tdata,
    input m_axis_fifo_118_tready,
    output ap_fifo_oarg_118_full_n,
    input [C_OUTPUT_FIFO_118_WIDTH-1:0] ap_fifo_oarg_118_din,
    input ap_fifo_oarg_118_write,
    //output FIFO to AXI-Stream interface 119
    output m_axis_fifo_119_tlast,
    output m_axis_fifo_119_tvalid,
    output [C_OUTPUT_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tkeep,
    output [C_OUTPUT_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tstrb,
    output [C_OUTPUT_FIFO_119_DMWIDTH-1:0] m_axis_fifo_119_tdata,
    input m_axis_fifo_119_tready,
    output ap_fifo_oarg_119_full_n,
    input [C_OUTPUT_FIFO_119_WIDTH-1:0] ap_fifo_oarg_119_din,
    input ap_fifo_oarg_119_write,
    //output FIFO to AXI-Stream interface 120
    output m_axis_fifo_120_tlast,
    output m_axis_fifo_120_tvalid,
    output [C_OUTPUT_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tkeep,
    output [C_OUTPUT_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tstrb,
    output [C_OUTPUT_FIFO_120_DMWIDTH-1:0] m_axis_fifo_120_tdata,
    input m_axis_fifo_120_tready,
    output ap_fifo_oarg_120_full_n,
    input [C_OUTPUT_FIFO_120_WIDTH-1:0] ap_fifo_oarg_120_din,
    input ap_fifo_oarg_120_write,
    //output FIFO to AXI-Stream interface 121
    output m_axis_fifo_121_tlast,
    output m_axis_fifo_121_tvalid,
    output [C_OUTPUT_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tkeep,
    output [C_OUTPUT_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tstrb,
    output [C_OUTPUT_FIFO_121_DMWIDTH-1:0] m_axis_fifo_121_tdata,
    input m_axis_fifo_121_tready,
    output ap_fifo_oarg_121_full_n,
    input [C_OUTPUT_FIFO_121_WIDTH-1:0] ap_fifo_oarg_121_din,
    input ap_fifo_oarg_121_write,
    //output FIFO to AXI-Stream interface 122
    output m_axis_fifo_122_tlast,
    output m_axis_fifo_122_tvalid,
    output [C_OUTPUT_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tkeep,
    output [C_OUTPUT_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tstrb,
    output [C_OUTPUT_FIFO_122_DMWIDTH-1:0] m_axis_fifo_122_tdata,
    input m_axis_fifo_122_tready,
    output ap_fifo_oarg_122_full_n,
    input [C_OUTPUT_FIFO_122_WIDTH-1:0] ap_fifo_oarg_122_din,
    input ap_fifo_oarg_122_write,
    //output FIFO to AXI-Stream interface 123
    output m_axis_fifo_123_tlast,
    output m_axis_fifo_123_tvalid,
    output [C_OUTPUT_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tkeep,
    output [C_OUTPUT_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tstrb,
    output [C_OUTPUT_FIFO_123_DMWIDTH-1:0] m_axis_fifo_123_tdata,
    input m_axis_fifo_123_tready,
    output ap_fifo_oarg_123_full_n,
    input [C_OUTPUT_FIFO_123_WIDTH-1:0] ap_fifo_oarg_123_din,
    input ap_fifo_oarg_123_write,
    //output FIFO to AXI-Stream interface 124
    output m_axis_fifo_124_tlast,
    output m_axis_fifo_124_tvalid,
    output [C_OUTPUT_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tkeep,
    output [C_OUTPUT_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tstrb,
    output [C_OUTPUT_FIFO_124_DMWIDTH-1:0] m_axis_fifo_124_tdata,
    input m_axis_fifo_124_tready,
    output ap_fifo_oarg_124_full_n,
    input [C_OUTPUT_FIFO_124_WIDTH-1:0] ap_fifo_oarg_124_din,
    input ap_fifo_oarg_124_write,
    //output FIFO to AXI-Stream interface 125
    output m_axis_fifo_125_tlast,
    output m_axis_fifo_125_tvalid,
    output [C_OUTPUT_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tkeep,
    output [C_OUTPUT_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tstrb,
    output [C_OUTPUT_FIFO_125_DMWIDTH-1:0] m_axis_fifo_125_tdata,
    input m_axis_fifo_125_tready,
    output ap_fifo_oarg_125_full_n,
    input [C_OUTPUT_FIFO_125_WIDTH-1:0] ap_fifo_oarg_125_din,
    input ap_fifo_oarg_125_write,
    //output FIFO to AXI-Stream interface 126
    output m_axis_fifo_126_tlast,
    output m_axis_fifo_126_tvalid,
    output [C_OUTPUT_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tkeep,
    output [C_OUTPUT_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tstrb,
    output [C_OUTPUT_FIFO_126_DMWIDTH-1:0] m_axis_fifo_126_tdata,
    input m_axis_fifo_126_tready,
    output ap_fifo_oarg_126_full_n,
    input [C_OUTPUT_FIFO_126_WIDTH-1:0] ap_fifo_oarg_126_din,
    input ap_fifo_oarg_126_write,
    //output FIFO to AXI-Stream interface 127
    output m_axis_fifo_127_tlast,
    output m_axis_fifo_127_tvalid,
    output [C_OUTPUT_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tkeep,
    output [C_OUTPUT_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tstrb,
    output [C_OUTPUT_FIFO_127_DMWIDTH-1:0] m_axis_fifo_127_tdata,
    input m_axis_fifo_127_tready,
    output ap_fifo_oarg_127_full_n,
    input [C_OUTPUT_FIFO_127_WIDTH-1:0] ap_fifo_oarg_127_din,
    input ap_fifo_oarg_127_write
    );

parameter C_NUM_OUTPUT_FIFOs = 0;
parameter [31:0] C_OUTPUT_FIFO_0_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_1_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_2_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_3_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_4_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_5_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_6_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_7_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_8_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_9_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_10_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_11_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_12_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_13_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_14_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_15_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_16_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_17_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_18_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_19_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_20_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_21_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_22_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_23_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_24_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_25_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_26_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_27_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_28_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_29_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_30_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_31_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_32_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_33_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_34_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_35_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_36_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_37_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_38_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_39_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_40_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_41_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_42_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_43_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_44_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_45_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_46_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_47_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_48_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_49_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_50_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_51_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_52_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_53_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_54_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_55_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_56_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_57_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_58_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_59_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_60_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_61_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_62_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_63_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_64_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_65_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_66_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_67_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_68_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_69_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_70_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_71_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_72_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_73_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_74_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_75_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_76_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_77_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_78_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_79_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_80_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_81_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_82_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_83_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_84_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_85_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_86_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_87_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_88_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_89_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_90_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_91_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_92_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_93_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_94_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_95_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_96_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_97_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_98_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_99_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_100_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_101_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_102_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_103_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_104_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_105_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_106_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_107_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_108_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_109_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_110_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_111_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_112_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_113_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_114_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_115_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_116_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_117_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_118_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_119_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_120_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_121_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_122_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_123_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_124_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_125_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_126_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_127_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_0_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_1_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_2_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_3_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_4_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_5_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_6_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_7_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_8_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_9_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_10_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_11_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_12_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_13_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_14_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_15_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_16_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_17_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_18_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_19_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_20_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_21_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_22_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_23_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_24_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_25_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_26_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_27_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_28_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_29_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_30_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_31_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_32_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_33_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_34_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_35_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_36_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_37_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_38_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_39_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_40_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_41_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_42_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_43_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_44_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_45_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_46_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_47_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_48_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_49_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_50_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_51_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_52_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_53_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_54_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_55_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_56_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_57_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_58_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_59_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_60_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_61_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_62_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_63_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_64_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_65_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_66_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_67_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_68_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_69_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_70_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_71_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_72_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_73_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_74_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_75_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_76_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_77_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_78_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_79_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_80_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_81_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_82_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_83_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_84_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_85_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_86_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_87_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_88_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_89_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_90_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_91_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_92_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_93_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_94_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_95_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_96_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_97_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_98_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_99_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_100_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_101_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_102_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_103_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_104_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_105_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_106_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_107_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_108_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_109_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_110_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_111_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_112_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_113_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_114_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_115_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_116_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_117_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_118_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_119_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_120_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_121_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_122_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_123_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_124_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_125_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_126_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_127_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_0_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_1_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_2_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_3_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_4_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_5_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_6_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_7_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_8_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_9_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_10_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_11_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_12_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_13_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_14_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_15_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_16_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_17_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_18_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_19_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_20_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_21_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_22_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_23_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_24_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_25_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_26_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_27_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_28_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_29_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_30_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_31_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_32_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_33_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_34_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_35_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_36_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_37_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_38_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_39_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_40_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_41_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_42_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_43_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_44_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_45_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_46_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_47_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_48_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_49_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_50_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_51_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_52_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_53_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_54_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_55_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_56_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_57_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_58_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_59_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_60_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_61_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_62_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_63_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_64_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_65_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_66_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_67_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_68_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_69_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_70_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_71_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_72_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_73_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_74_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_75_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_76_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_77_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_78_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_79_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_80_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_81_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_82_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_83_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_84_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_85_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_86_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_87_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_88_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_89_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_90_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_91_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_92_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_93_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_94_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_95_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_96_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_97_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_98_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_99_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_100_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_101_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_102_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_103_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_104_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_105_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_106_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_107_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_108_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_109_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_110_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_111_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_112_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_113_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_114_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_115_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_116_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_117_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_118_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_119_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_120_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_121_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_122_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_123_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_124_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_125_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_126_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_127_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface

    localparam C_MAX_OUTPUT_FIFOs = 128;
    localparam C_MAX_BIT_WIDTH = 1024;
    localparam [(C_MAX_OUTPUT_FIFOs*32)-1:0] C_OUTFIFO_BIT_ARRAY = {C_OUTPUT_FIFO_127_WIDTH,C_OUTPUT_FIFO_126_WIDTH,C_OUTPUT_FIFO_125_WIDTH,C_OUTPUT_FIFO_124_WIDTH,C_OUTPUT_FIFO_123_WIDTH,C_OUTPUT_FIFO_122_WIDTH,C_OUTPUT_FIFO_121_WIDTH,C_OUTPUT_FIFO_120_WIDTH,C_OUTPUT_FIFO_119_WIDTH,C_OUTPUT_FIFO_118_WIDTH,C_OUTPUT_FIFO_117_WIDTH,C_OUTPUT_FIFO_116_WIDTH,C_OUTPUT_FIFO_115_WIDTH,C_OUTPUT_FIFO_114_WIDTH,C_OUTPUT_FIFO_113_WIDTH,C_OUTPUT_FIFO_112_WIDTH,C_OUTPUT_FIFO_111_WIDTH,C_OUTPUT_FIFO_110_WIDTH,C_OUTPUT_FIFO_109_WIDTH,C_OUTPUT_FIFO_108_WIDTH,C_OUTPUT_FIFO_107_WIDTH,C_OUTPUT_FIFO_106_WIDTH,C_OUTPUT_FIFO_105_WIDTH,C_OUTPUT_FIFO_104_WIDTH,C_OUTPUT_FIFO_103_WIDTH,C_OUTPUT_FIFO_102_WIDTH,C_OUTPUT_FIFO_101_WIDTH,C_OUTPUT_FIFO_100_WIDTH,C_OUTPUT_FIFO_99_WIDTH,C_OUTPUT_FIFO_98_WIDTH,C_OUTPUT_FIFO_97_WIDTH,C_OUTPUT_FIFO_96_WIDTH,C_OUTPUT_FIFO_95_WIDTH,C_OUTPUT_FIFO_94_WIDTH,C_OUTPUT_FIFO_93_WIDTH,C_OUTPUT_FIFO_92_WIDTH,C_OUTPUT_FIFO_91_WIDTH,C_OUTPUT_FIFO_90_WIDTH,C_OUTPUT_FIFO_89_WIDTH,C_OUTPUT_FIFO_88_WIDTH,C_OUTPUT_FIFO_87_WIDTH,C_OUTPUT_FIFO_86_WIDTH,C_OUTPUT_FIFO_85_WIDTH,C_OUTPUT_FIFO_84_WIDTH,C_OUTPUT_FIFO_83_WIDTH,C_OUTPUT_FIFO_82_WIDTH,C_OUTPUT_FIFO_81_WIDTH,C_OUTPUT_FIFO_80_WIDTH,C_OUTPUT_FIFO_79_WIDTH,C_OUTPUT_FIFO_78_WIDTH,C_OUTPUT_FIFO_77_WIDTH,C_OUTPUT_FIFO_76_WIDTH,C_OUTPUT_FIFO_75_WIDTH,C_OUTPUT_FIFO_74_WIDTH,C_OUTPUT_FIFO_73_WIDTH,C_OUTPUT_FIFO_72_WIDTH,C_OUTPUT_FIFO_71_WIDTH,C_OUTPUT_FIFO_70_WIDTH,C_OUTPUT_FIFO_69_WIDTH,C_OUTPUT_FIFO_68_WIDTH,C_OUTPUT_FIFO_67_WIDTH,C_OUTPUT_FIFO_66_WIDTH,C_OUTPUT_FIFO_65_WIDTH,C_OUTPUT_FIFO_64_WIDTH,C_OUTPUT_FIFO_63_WIDTH,C_OUTPUT_FIFO_62_WIDTH,C_OUTPUT_FIFO_61_WIDTH,C_OUTPUT_FIFO_60_WIDTH,C_OUTPUT_FIFO_59_WIDTH,C_OUTPUT_FIFO_58_WIDTH,C_OUTPUT_FIFO_57_WIDTH,C_OUTPUT_FIFO_56_WIDTH,C_OUTPUT_FIFO_55_WIDTH,C_OUTPUT_FIFO_54_WIDTH,C_OUTPUT_FIFO_53_WIDTH,C_OUTPUT_FIFO_52_WIDTH,C_OUTPUT_FIFO_51_WIDTH,C_OUTPUT_FIFO_50_WIDTH,C_OUTPUT_FIFO_49_WIDTH,C_OUTPUT_FIFO_48_WIDTH,C_OUTPUT_FIFO_47_WIDTH,C_OUTPUT_FIFO_46_WIDTH,C_OUTPUT_FIFO_45_WIDTH,C_OUTPUT_FIFO_44_WIDTH,C_OUTPUT_FIFO_43_WIDTH,C_OUTPUT_FIFO_42_WIDTH,C_OUTPUT_FIFO_41_WIDTH,C_OUTPUT_FIFO_40_WIDTH,C_OUTPUT_FIFO_39_WIDTH,C_OUTPUT_FIFO_38_WIDTH,C_OUTPUT_FIFO_37_WIDTH,C_OUTPUT_FIFO_36_WIDTH,C_OUTPUT_FIFO_35_WIDTH,C_OUTPUT_FIFO_34_WIDTH,C_OUTPUT_FIFO_33_WIDTH,C_OUTPUT_FIFO_32_WIDTH,C_OUTPUT_FIFO_31_WIDTH,C_OUTPUT_FIFO_30_WIDTH,C_OUTPUT_FIFO_29_WIDTH,C_OUTPUT_FIFO_28_WIDTH,C_OUTPUT_FIFO_27_WIDTH,C_OUTPUT_FIFO_26_WIDTH,C_OUTPUT_FIFO_25_WIDTH,C_OUTPUT_FIFO_24_WIDTH,C_OUTPUT_FIFO_23_WIDTH,C_OUTPUT_FIFO_22_WIDTH,C_OUTPUT_FIFO_21_WIDTH,C_OUTPUT_FIFO_20_WIDTH,C_OUTPUT_FIFO_19_WIDTH,C_OUTPUT_FIFO_18_WIDTH,C_OUTPUT_FIFO_17_WIDTH,C_OUTPUT_FIFO_16_WIDTH,C_OUTPUT_FIFO_15_WIDTH,C_OUTPUT_FIFO_14_WIDTH,C_OUTPUT_FIFO_13_WIDTH,C_OUTPUT_FIFO_12_WIDTH,C_OUTPUT_FIFO_11_WIDTH,C_OUTPUT_FIFO_10_WIDTH,C_OUTPUT_FIFO_9_WIDTH,C_OUTPUT_FIFO_8_WIDTH,C_OUTPUT_FIFO_7_WIDTH,C_OUTPUT_FIFO_6_WIDTH,C_OUTPUT_FIFO_5_WIDTH,C_OUTPUT_FIFO_4_WIDTH,C_OUTPUT_FIFO_3_WIDTH,C_OUTPUT_FIFO_2_WIDTH,C_OUTPUT_FIFO_1_WIDTH,C_OUTPUT_FIFO_0_WIDTH};
    localparam [(C_MAX_OUTPUT_FIFOs*32)-1:0] C_DEPTH_BIT_ARRAY = {C_OUTPUT_FIFO_127_DEPTH,C_OUTPUT_FIFO_126_DEPTH,C_OUTPUT_FIFO_125_DEPTH,C_OUTPUT_FIFO_124_DEPTH,C_OUTPUT_FIFO_123_DEPTH,C_OUTPUT_FIFO_122_DEPTH,C_OUTPUT_FIFO_121_DEPTH,C_OUTPUT_FIFO_120_DEPTH,C_OUTPUT_FIFO_119_DEPTH,C_OUTPUT_FIFO_118_DEPTH,C_OUTPUT_FIFO_117_DEPTH,C_OUTPUT_FIFO_116_DEPTH,C_OUTPUT_FIFO_115_DEPTH,C_OUTPUT_FIFO_114_DEPTH,C_OUTPUT_FIFO_113_DEPTH,C_OUTPUT_FIFO_112_DEPTH,C_OUTPUT_FIFO_111_DEPTH,C_OUTPUT_FIFO_110_DEPTH,C_OUTPUT_FIFO_109_DEPTH,C_OUTPUT_FIFO_108_DEPTH,C_OUTPUT_FIFO_107_DEPTH,C_OUTPUT_FIFO_106_DEPTH,C_OUTPUT_FIFO_105_DEPTH,C_OUTPUT_FIFO_104_DEPTH,C_OUTPUT_FIFO_103_DEPTH,C_OUTPUT_FIFO_102_DEPTH,C_OUTPUT_FIFO_101_DEPTH,C_OUTPUT_FIFO_100_DEPTH,C_OUTPUT_FIFO_99_DEPTH,C_OUTPUT_FIFO_98_DEPTH,C_OUTPUT_FIFO_97_DEPTH,C_OUTPUT_FIFO_96_DEPTH,C_OUTPUT_FIFO_95_DEPTH,C_OUTPUT_FIFO_94_DEPTH,C_OUTPUT_FIFO_93_DEPTH,C_OUTPUT_FIFO_92_DEPTH,C_OUTPUT_FIFO_91_DEPTH,C_OUTPUT_FIFO_90_DEPTH,C_OUTPUT_FIFO_89_DEPTH,C_OUTPUT_FIFO_88_DEPTH,C_OUTPUT_FIFO_87_DEPTH,C_OUTPUT_FIFO_86_DEPTH,C_OUTPUT_FIFO_85_DEPTH,C_OUTPUT_FIFO_84_DEPTH,C_OUTPUT_FIFO_83_DEPTH,C_OUTPUT_FIFO_82_DEPTH,C_OUTPUT_FIFO_81_DEPTH,C_OUTPUT_FIFO_80_DEPTH,C_OUTPUT_FIFO_79_DEPTH,C_OUTPUT_FIFO_78_DEPTH,C_OUTPUT_FIFO_77_DEPTH,C_OUTPUT_FIFO_76_DEPTH,C_OUTPUT_FIFO_75_DEPTH,C_OUTPUT_FIFO_74_DEPTH,C_OUTPUT_FIFO_73_DEPTH,C_OUTPUT_FIFO_72_DEPTH,C_OUTPUT_FIFO_71_DEPTH,C_OUTPUT_FIFO_70_DEPTH,C_OUTPUT_FIFO_69_DEPTH,C_OUTPUT_FIFO_68_DEPTH,C_OUTPUT_FIFO_67_DEPTH,C_OUTPUT_FIFO_66_DEPTH,C_OUTPUT_FIFO_65_DEPTH,C_OUTPUT_FIFO_64_DEPTH,C_OUTPUT_FIFO_63_DEPTH,C_OUTPUT_FIFO_62_DEPTH,C_OUTPUT_FIFO_61_DEPTH,C_OUTPUT_FIFO_60_DEPTH,C_OUTPUT_FIFO_59_DEPTH,C_OUTPUT_FIFO_58_DEPTH,C_OUTPUT_FIFO_57_DEPTH,C_OUTPUT_FIFO_56_DEPTH,C_OUTPUT_FIFO_55_DEPTH,C_OUTPUT_FIFO_54_DEPTH,C_OUTPUT_FIFO_53_DEPTH,C_OUTPUT_FIFO_52_DEPTH,C_OUTPUT_FIFO_51_DEPTH,C_OUTPUT_FIFO_50_DEPTH,C_OUTPUT_FIFO_49_DEPTH,C_OUTPUT_FIFO_48_DEPTH,C_OUTPUT_FIFO_47_DEPTH,C_OUTPUT_FIFO_46_DEPTH,C_OUTPUT_FIFO_45_DEPTH,C_OUTPUT_FIFO_44_DEPTH,C_OUTPUT_FIFO_43_DEPTH,C_OUTPUT_FIFO_42_DEPTH,C_OUTPUT_FIFO_41_DEPTH,C_OUTPUT_FIFO_40_DEPTH,C_OUTPUT_FIFO_39_DEPTH,C_OUTPUT_FIFO_38_DEPTH,C_OUTPUT_FIFO_37_DEPTH,C_OUTPUT_FIFO_36_DEPTH,C_OUTPUT_FIFO_35_DEPTH,C_OUTPUT_FIFO_34_DEPTH,C_OUTPUT_FIFO_33_DEPTH,C_OUTPUT_FIFO_32_DEPTH,C_OUTPUT_FIFO_31_DEPTH,C_OUTPUT_FIFO_30_DEPTH,C_OUTPUT_FIFO_29_DEPTH,C_OUTPUT_FIFO_28_DEPTH,C_OUTPUT_FIFO_27_DEPTH,C_OUTPUT_FIFO_26_DEPTH,C_OUTPUT_FIFO_25_DEPTH,C_OUTPUT_FIFO_24_DEPTH,C_OUTPUT_FIFO_23_DEPTH,C_OUTPUT_FIFO_22_DEPTH,C_OUTPUT_FIFO_21_DEPTH,C_OUTPUT_FIFO_20_DEPTH,C_OUTPUT_FIFO_19_DEPTH,C_OUTPUT_FIFO_18_DEPTH,C_OUTPUT_FIFO_17_DEPTH,C_OUTPUT_FIFO_16_DEPTH,C_OUTPUT_FIFO_15_DEPTH,C_OUTPUT_FIFO_14_DEPTH,C_OUTPUT_FIFO_13_DEPTH,C_OUTPUT_FIFO_12_DEPTH,C_OUTPUT_FIFO_11_DEPTH,C_OUTPUT_FIFO_10_DEPTH,C_OUTPUT_FIFO_9_DEPTH,C_OUTPUT_FIFO_8_DEPTH,C_OUTPUT_FIFO_7_DEPTH,C_OUTPUT_FIFO_6_DEPTH,C_OUTPUT_FIFO_5_DEPTH,C_OUTPUT_FIFO_4_DEPTH,C_OUTPUT_FIFO_3_DEPTH,C_OUTPUT_FIFO_2_DEPTH,C_OUTPUT_FIFO_1_DEPTH,C_OUTPUT_FIFO_0_DEPTH};
    localparam [(C_MAX_OUTPUT_FIFOs*32)-1:0] C_DMWIDTH_BIT_ARRAY = {C_OUTPUT_FIFO_127_DMWIDTH,C_OUTPUT_FIFO_126_DMWIDTH,C_OUTPUT_FIFO_125_DMWIDTH,C_OUTPUT_FIFO_124_DMWIDTH,C_OUTPUT_FIFO_123_DMWIDTH,C_OUTPUT_FIFO_122_DMWIDTH,C_OUTPUT_FIFO_121_DMWIDTH,C_OUTPUT_FIFO_120_DMWIDTH,C_OUTPUT_FIFO_119_DMWIDTH,C_OUTPUT_FIFO_118_DMWIDTH,C_OUTPUT_FIFO_117_DMWIDTH,C_OUTPUT_FIFO_116_DMWIDTH,C_OUTPUT_FIFO_115_DMWIDTH,C_OUTPUT_FIFO_114_DMWIDTH,C_OUTPUT_FIFO_113_DMWIDTH,C_OUTPUT_FIFO_112_DMWIDTH,C_OUTPUT_FIFO_111_DMWIDTH,C_OUTPUT_FIFO_110_DMWIDTH,C_OUTPUT_FIFO_109_DMWIDTH,C_OUTPUT_FIFO_108_DMWIDTH,C_OUTPUT_FIFO_107_DMWIDTH,C_OUTPUT_FIFO_106_DMWIDTH,C_OUTPUT_FIFO_105_DMWIDTH,C_OUTPUT_FIFO_104_DMWIDTH,C_OUTPUT_FIFO_103_DMWIDTH,C_OUTPUT_FIFO_102_DMWIDTH,C_OUTPUT_FIFO_101_DMWIDTH,C_OUTPUT_FIFO_100_DMWIDTH,C_OUTPUT_FIFO_99_DMWIDTH,C_OUTPUT_FIFO_98_DMWIDTH,C_OUTPUT_FIFO_97_DMWIDTH,C_OUTPUT_FIFO_96_DMWIDTH,C_OUTPUT_FIFO_95_DMWIDTH,C_OUTPUT_FIFO_94_DMWIDTH,C_OUTPUT_FIFO_93_DMWIDTH,C_OUTPUT_FIFO_92_DMWIDTH,C_OUTPUT_FIFO_91_DMWIDTH,C_OUTPUT_FIFO_90_DMWIDTH,C_OUTPUT_FIFO_89_DMWIDTH,C_OUTPUT_FIFO_88_DMWIDTH,C_OUTPUT_FIFO_87_DMWIDTH,C_OUTPUT_FIFO_86_DMWIDTH,C_OUTPUT_FIFO_85_DMWIDTH,C_OUTPUT_FIFO_84_DMWIDTH,C_OUTPUT_FIFO_83_DMWIDTH,C_OUTPUT_FIFO_82_DMWIDTH,C_OUTPUT_FIFO_81_DMWIDTH,C_OUTPUT_FIFO_80_DMWIDTH,C_OUTPUT_FIFO_79_DMWIDTH,C_OUTPUT_FIFO_78_DMWIDTH,C_OUTPUT_FIFO_77_DMWIDTH,C_OUTPUT_FIFO_76_DMWIDTH,C_OUTPUT_FIFO_75_DMWIDTH,C_OUTPUT_FIFO_74_DMWIDTH,C_OUTPUT_FIFO_73_DMWIDTH,C_OUTPUT_FIFO_72_DMWIDTH,C_OUTPUT_FIFO_71_DMWIDTH,C_OUTPUT_FIFO_70_DMWIDTH,C_OUTPUT_FIFO_69_DMWIDTH,C_OUTPUT_FIFO_68_DMWIDTH,C_OUTPUT_FIFO_67_DMWIDTH,C_OUTPUT_FIFO_66_DMWIDTH,C_OUTPUT_FIFO_65_DMWIDTH,C_OUTPUT_FIFO_64_DMWIDTH,C_OUTPUT_FIFO_63_DMWIDTH,C_OUTPUT_FIFO_62_DMWIDTH,C_OUTPUT_FIFO_61_DMWIDTH,C_OUTPUT_FIFO_60_DMWIDTH,C_OUTPUT_FIFO_59_DMWIDTH,C_OUTPUT_FIFO_58_DMWIDTH,C_OUTPUT_FIFO_57_DMWIDTH,C_OUTPUT_FIFO_56_DMWIDTH,C_OUTPUT_FIFO_55_DMWIDTH,C_OUTPUT_FIFO_54_DMWIDTH,C_OUTPUT_FIFO_53_DMWIDTH,C_OUTPUT_FIFO_52_DMWIDTH,C_OUTPUT_FIFO_51_DMWIDTH,C_OUTPUT_FIFO_50_DMWIDTH,C_OUTPUT_FIFO_49_DMWIDTH,C_OUTPUT_FIFO_48_DMWIDTH,C_OUTPUT_FIFO_47_DMWIDTH,C_OUTPUT_FIFO_46_DMWIDTH,C_OUTPUT_FIFO_45_DMWIDTH,C_OUTPUT_FIFO_44_DMWIDTH,C_OUTPUT_FIFO_43_DMWIDTH,C_OUTPUT_FIFO_42_DMWIDTH,C_OUTPUT_FIFO_41_DMWIDTH,C_OUTPUT_FIFO_40_DMWIDTH,C_OUTPUT_FIFO_39_DMWIDTH,C_OUTPUT_FIFO_38_DMWIDTH,C_OUTPUT_FIFO_37_DMWIDTH,C_OUTPUT_FIFO_36_DMWIDTH,C_OUTPUT_FIFO_35_DMWIDTH,C_OUTPUT_FIFO_34_DMWIDTH,C_OUTPUT_FIFO_33_DMWIDTH,C_OUTPUT_FIFO_32_DMWIDTH,C_OUTPUT_FIFO_31_DMWIDTH,C_OUTPUT_FIFO_30_DMWIDTH,C_OUTPUT_FIFO_29_DMWIDTH,C_OUTPUT_FIFO_28_DMWIDTH,C_OUTPUT_FIFO_27_DMWIDTH,C_OUTPUT_FIFO_26_DMWIDTH,C_OUTPUT_FIFO_25_DMWIDTH,C_OUTPUT_FIFO_24_DMWIDTH,C_OUTPUT_FIFO_23_DMWIDTH,C_OUTPUT_FIFO_22_DMWIDTH,C_OUTPUT_FIFO_21_DMWIDTH,C_OUTPUT_FIFO_20_DMWIDTH,C_OUTPUT_FIFO_19_DMWIDTH,C_OUTPUT_FIFO_18_DMWIDTH,C_OUTPUT_FIFO_17_DMWIDTH,C_OUTPUT_FIFO_16_DMWIDTH,C_OUTPUT_FIFO_15_DMWIDTH,C_OUTPUT_FIFO_14_DMWIDTH,C_OUTPUT_FIFO_13_DMWIDTH,C_OUTPUT_FIFO_12_DMWIDTH,C_OUTPUT_FIFO_11_DMWIDTH,C_OUTPUT_FIFO_10_DMWIDTH,C_OUTPUT_FIFO_9_DMWIDTH,C_OUTPUT_FIFO_8_DMWIDTH,C_OUTPUT_FIFO_7_DMWIDTH,C_OUTPUT_FIFO_6_DMWIDTH,C_OUTPUT_FIFO_5_DMWIDTH,C_OUTPUT_FIFO_4_DMWIDTH,C_OUTPUT_FIFO_3_DMWIDTH,C_OUTPUT_FIFO_2_DMWIDTH,C_OUTPUT_FIFO_1_DMWIDTH,C_OUTPUT_FIFO_0_DMWIDTH};
    
    wire [C_MAX_OUTPUT_FIFOs-1:0] tlast;
    wire [C_MAX_OUTPUT_FIFOs-1:0] tvalid;
    wire [C_MAX_OUTPUT_FIFOs-1:0] tready;
    wire [C_MAX_BIT_WIDTH/8-1:0] tkeep [C_NUM_OUTPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] tstrb [C_NUM_OUTPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0] tdata [C_MAX_OUTPUT_FIFOs-1:0];
    
    wire [C_MAX_OUTPUT_FIFOs-1:0] buf_tlast;
    wire [C_MAX_OUTPUT_FIFOs-1:0] buf_tvalid;
    wire [C_MAX_OUTPUT_FIFOs-1:0] buf_tready;
    wire [C_MAX_BIT_WIDTH-1:0] buf_tdata [C_MAX_OUTPUT_FIFOs-1:0];
    
    wire [C_MAX_OUTPUT_FIFOs-1:0] dwconv_tlast;
    wire [C_MAX_OUTPUT_FIFOs-1:0] dwconv_tvalid;
    wire [C_MAX_OUTPUT_FIFOs-1:0] dwconv_tready;
    wire [C_MAX_BIT_WIDTH/8-1:0] dwconv_tkeep [C_NUM_OUTPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] dwconv_tstrb [C_NUM_OUTPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0] dwconv_tdata [C_MAX_OUTPUT_FIFOs-1:0];
    
    wire [C_MAX_OUTPUT_FIFOs-1:0] write;
    wire [C_MAX_OUTPUT_FIFOs-1:0] full;
    wire [C_MAX_BIT_WIDTH-1:0] din [C_MAX_OUTPUT_FIFOs-1:0];
        
    //assign inputs to buses, and buses to outputs
    generate
        if(C_NUM_OUTPUT_FIFOs > 0) begin
            assign dwconv_tready[0] = m_axis_fifo_0_tready;
            assign m_axis_fifo_0_tlast = dwconv_tlast[0];
            assign m_axis_fifo_0_tvalid = dwconv_tvalid[0];
            assign m_axis_fifo_0_tkeep = dwconv_tkeep[0][C_OUTPUT_FIFO_0_DMWIDTH/8-1:0];
            assign m_axis_fifo_0_tstrb = dwconv_tstrb[0][C_OUTPUT_FIFO_0_DMWIDTH/8-1:0];
            assign m_axis_fifo_0_tdata = dwconv_tdata[0][C_OUTPUT_FIFO_0_DMWIDTH-1:0];
            assign ap_fifo_oarg_0_full_n = full[0];
            assign write[0] = ap_fifo_oarg_0_write;
            assign din[0][C_OUTPUT_FIFO_0_WIDTH-1:0] = ap_fifo_oarg_0_din;
            assign tkeep[0] = {C_OUTPUT_FIFO_0_WIDTH/8{1'b1}};
            assign tstrb[0] = {C_OUTPUT_FIFO_0_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 1) begin
            assign dwconv_tready[1] = m_axis_fifo_1_tready;
            assign m_axis_fifo_1_tlast = dwconv_tlast[1];
            assign m_axis_fifo_1_tvalid = dwconv_tvalid[1];
            assign m_axis_fifo_1_tkeep = dwconv_tkeep[1][C_OUTPUT_FIFO_1_DMWIDTH/8-1:0];
            assign m_axis_fifo_1_tstrb = dwconv_tstrb[1][C_OUTPUT_FIFO_1_DMWIDTH/8-1:0];
            assign m_axis_fifo_1_tdata = dwconv_tdata[1][C_OUTPUT_FIFO_1_DMWIDTH-1:0];
            assign ap_fifo_oarg_1_full_n = full[1];
            assign write[1] = ap_fifo_oarg_1_write;
            assign din[1][C_OUTPUT_FIFO_1_WIDTH-1:0] = ap_fifo_oarg_1_din;
            assign tkeep[1] = {C_OUTPUT_FIFO_1_WIDTH/8{1'b1}};
            assign tstrb[1] = {C_OUTPUT_FIFO_1_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 2) begin
            assign dwconv_tready[2] = m_axis_fifo_2_tready;
            assign m_axis_fifo_2_tlast = dwconv_tlast[2];
            assign m_axis_fifo_2_tvalid = dwconv_tvalid[2];
            assign m_axis_fifo_2_tkeep = dwconv_tkeep[2][C_OUTPUT_FIFO_2_DMWIDTH/8-1:0];
            assign m_axis_fifo_2_tstrb = dwconv_tstrb[2][C_OUTPUT_FIFO_2_DMWIDTH/8-1:0];
            assign m_axis_fifo_2_tdata = dwconv_tdata[2][C_OUTPUT_FIFO_2_DMWIDTH-1:0];
            assign ap_fifo_oarg_2_full_n = full[2];
            assign write[2] = ap_fifo_oarg_2_write;
            assign din[2][C_OUTPUT_FIFO_2_WIDTH-1:0] = ap_fifo_oarg_2_din;
            assign tkeep[2] = {C_OUTPUT_FIFO_2_WIDTH/8{1'b1}};
            assign tstrb[2] = {C_OUTPUT_FIFO_2_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 3) begin
            assign dwconv_tready[3] = m_axis_fifo_3_tready;
            assign m_axis_fifo_3_tlast = dwconv_tlast[3];
            assign m_axis_fifo_3_tvalid = dwconv_tvalid[3];
            assign m_axis_fifo_3_tkeep = dwconv_tkeep[3][C_OUTPUT_FIFO_3_DMWIDTH/8-1:0];
            assign m_axis_fifo_3_tstrb = dwconv_tstrb[3][C_OUTPUT_FIFO_3_DMWIDTH/8-1:0];
            assign m_axis_fifo_3_tdata = dwconv_tdata[3][C_OUTPUT_FIFO_3_DMWIDTH-1:0];
            assign ap_fifo_oarg_3_full_n = full[3];
            assign write[3] = ap_fifo_oarg_3_write;
            assign din[3][C_OUTPUT_FIFO_3_WIDTH-1:0] = ap_fifo_oarg_3_din;
            assign tkeep[3] = {C_OUTPUT_FIFO_3_WIDTH/8{1'b1}};
            assign tstrb[3] = {C_OUTPUT_FIFO_3_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 4) begin
            assign dwconv_tready[4] = m_axis_fifo_4_tready;
            assign m_axis_fifo_4_tlast = dwconv_tlast[4];
            assign m_axis_fifo_4_tvalid = dwconv_tvalid[4];
            assign m_axis_fifo_4_tkeep = dwconv_tkeep[4][C_OUTPUT_FIFO_4_DMWIDTH/8-1:0];
            assign m_axis_fifo_4_tstrb = dwconv_tstrb[4][C_OUTPUT_FIFO_4_DMWIDTH/8-1:0];
            assign m_axis_fifo_4_tdata = dwconv_tdata[4][C_OUTPUT_FIFO_4_DMWIDTH-1:0];
            assign ap_fifo_oarg_4_full_n = full[4];
            assign write[4] = ap_fifo_oarg_4_write;
            assign din[4][C_OUTPUT_FIFO_4_WIDTH-1:0] = ap_fifo_oarg_4_din;
            assign tkeep[4] = {C_OUTPUT_FIFO_4_WIDTH/8{1'b1}};
            assign tstrb[4] = {C_OUTPUT_FIFO_4_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 5) begin
            assign dwconv_tready[5] = m_axis_fifo_5_tready;
            assign m_axis_fifo_5_tlast = dwconv_tlast[5];
            assign m_axis_fifo_5_tvalid = dwconv_tvalid[5];
            assign m_axis_fifo_5_tkeep = dwconv_tkeep[5][C_OUTPUT_FIFO_5_DMWIDTH/8-1:0];
            assign m_axis_fifo_5_tstrb = dwconv_tstrb[5][C_OUTPUT_FIFO_5_DMWIDTH/8-1:0];
            assign m_axis_fifo_5_tdata = dwconv_tdata[5][C_OUTPUT_FIFO_5_DMWIDTH-1:0];
            assign ap_fifo_oarg_5_full_n = full[5];
            assign write[5] = ap_fifo_oarg_5_write;
            assign din[5][C_OUTPUT_FIFO_5_WIDTH-1:0] = ap_fifo_oarg_5_din;
            assign tkeep[5] = {C_OUTPUT_FIFO_5_WIDTH/8{1'b1}};
            assign tstrb[5] = {C_OUTPUT_FIFO_5_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 6) begin
            assign dwconv_tready[6] = m_axis_fifo_6_tready;
            assign m_axis_fifo_6_tlast = dwconv_tlast[6];
            assign m_axis_fifo_6_tvalid = dwconv_tvalid[6];
            assign m_axis_fifo_6_tkeep = dwconv_tkeep[6][C_OUTPUT_FIFO_6_DMWIDTH/8-1:0];
            assign m_axis_fifo_6_tstrb = dwconv_tstrb[6][C_OUTPUT_FIFO_6_DMWIDTH/8-1:0];
            assign m_axis_fifo_6_tdata = dwconv_tdata[6][C_OUTPUT_FIFO_6_DMWIDTH-1:0];
            assign ap_fifo_oarg_6_full_n = full[6];
            assign write[6] = ap_fifo_oarg_6_write;
            assign din[6][C_OUTPUT_FIFO_6_WIDTH-1:0] = ap_fifo_oarg_6_din;
            assign tkeep[6] = {C_OUTPUT_FIFO_6_WIDTH/8{1'b1}};
            assign tstrb[6] = {C_OUTPUT_FIFO_6_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 7) begin
            assign dwconv_tready[7] = m_axis_fifo_7_tready;
            assign m_axis_fifo_7_tlast = dwconv_tlast[7];
            assign m_axis_fifo_7_tvalid = dwconv_tvalid[7];
            assign m_axis_fifo_7_tkeep = dwconv_tkeep[7][C_OUTPUT_FIFO_7_DMWIDTH/8-1:0];
            assign m_axis_fifo_7_tstrb = dwconv_tstrb[7][C_OUTPUT_FIFO_7_DMWIDTH/8-1:0];
            assign m_axis_fifo_7_tdata = dwconv_tdata[7][C_OUTPUT_FIFO_7_DMWIDTH-1:0];
            assign ap_fifo_oarg_7_full_n = full[7];
            assign write[7] = ap_fifo_oarg_7_write;
            assign din[7][C_OUTPUT_FIFO_7_WIDTH-1:0] = ap_fifo_oarg_7_din;
            assign tkeep[7] = {C_OUTPUT_FIFO_7_WIDTH/8{1'b1}};
            assign tstrb[7] = {C_OUTPUT_FIFO_7_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 8) begin
            assign dwconv_tready[8] = m_axis_fifo_8_tready;
            assign m_axis_fifo_8_tlast = dwconv_tlast[8];
            assign m_axis_fifo_8_tvalid = dwconv_tvalid[8];
            assign m_axis_fifo_8_tkeep = dwconv_tkeep[8][C_OUTPUT_FIFO_8_DMWIDTH/8-1:0];
            assign m_axis_fifo_8_tstrb = dwconv_tstrb[8][C_OUTPUT_FIFO_8_DMWIDTH/8-1:0];
            assign m_axis_fifo_8_tdata = dwconv_tdata[8][C_OUTPUT_FIFO_8_DMWIDTH-1:0];
            assign ap_fifo_oarg_8_full_n = full[8];
            assign write[8] = ap_fifo_oarg_8_write;
            assign din[8][C_OUTPUT_FIFO_8_WIDTH-1:0] = ap_fifo_oarg_8_din;
            assign tkeep[8] = {C_OUTPUT_FIFO_8_WIDTH/8{1'b1}};
            assign tstrb[8] = {C_OUTPUT_FIFO_8_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 9) begin
            assign dwconv_tready[9] = m_axis_fifo_9_tready;
            assign m_axis_fifo_9_tlast = dwconv_tlast[9];
            assign m_axis_fifo_9_tvalid = dwconv_tvalid[9];
            assign m_axis_fifo_9_tkeep = dwconv_tkeep[9][C_OUTPUT_FIFO_9_DMWIDTH/8-1:0];
            assign m_axis_fifo_9_tstrb = dwconv_tstrb[9][C_OUTPUT_FIFO_9_DMWIDTH/8-1:0];
            assign m_axis_fifo_9_tdata = dwconv_tdata[9][C_OUTPUT_FIFO_9_DMWIDTH-1:0];
            assign ap_fifo_oarg_9_full_n = full[9];
            assign write[9] = ap_fifo_oarg_9_write;
            assign din[9][C_OUTPUT_FIFO_9_WIDTH-1:0] = ap_fifo_oarg_9_din;
            assign tkeep[9] = {C_OUTPUT_FIFO_9_WIDTH/8{1'b1}};
            assign tstrb[9] = {C_OUTPUT_FIFO_9_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 10) begin
            assign dwconv_tready[10] = m_axis_fifo_10_tready;
            assign m_axis_fifo_10_tlast = dwconv_tlast[10];
            assign m_axis_fifo_10_tvalid = dwconv_tvalid[10];
            assign m_axis_fifo_10_tkeep = dwconv_tkeep[10][C_OUTPUT_FIFO_10_DMWIDTH/8-1:0];
            assign m_axis_fifo_10_tstrb = dwconv_tstrb[10][C_OUTPUT_FIFO_10_DMWIDTH/8-1:0];
            assign m_axis_fifo_10_tdata = dwconv_tdata[10][C_OUTPUT_FIFO_10_DMWIDTH-1:0];
            assign ap_fifo_oarg_10_full_n = full[10];
            assign write[10] = ap_fifo_oarg_10_write;
            assign din[10][C_OUTPUT_FIFO_10_WIDTH-1:0] = ap_fifo_oarg_10_din;
            assign tkeep[10] = {C_OUTPUT_FIFO_10_WIDTH/8{1'b1}};
            assign tstrb[10] = {C_OUTPUT_FIFO_10_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 11) begin
            assign dwconv_tready[11] = m_axis_fifo_11_tready;
            assign m_axis_fifo_11_tlast = dwconv_tlast[11];
            assign m_axis_fifo_11_tvalid = dwconv_tvalid[11];
            assign m_axis_fifo_11_tkeep = dwconv_tkeep[11][C_OUTPUT_FIFO_11_DMWIDTH/8-1:0];
            assign m_axis_fifo_11_tstrb = dwconv_tstrb[11][C_OUTPUT_FIFO_11_DMWIDTH/8-1:0];
            assign m_axis_fifo_11_tdata = dwconv_tdata[11][C_OUTPUT_FIFO_11_DMWIDTH-1:0];
            assign ap_fifo_oarg_11_full_n = full[11];
            assign write[11] = ap_fifo_oarg_11_write;
            assign din[11][C_OUTPUT_FIFO_11_WIDTH-1:0] = ap_fifo_oarg_11_din;
            assign tkeep[11] = {C_OUTPUT_FIFO_11_WIDTH/8{1'b1}};
            assign tstrb[11] = {C_OUTPUT_FIFO_11_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 12) begin
            assign dwconv_tready[12] = m_axis_fifo_12_tready;
            assign m_axis_fifo_12_tlast = dwconv_tlast[12];
            assign m_axis_fifo_12_tvalid = dwconv_tvalid[12];
            assign m_axis_fifo_12_tkeep = dwconv_tkeep[12][C_OUTPUT_FIFO_12_DMWIDTH/8-1:0];
            assign m_axis_fifo_12_tstrb = dwconv_tstrb[12][C_OUTPUT_FIFO_12_DMWIDTH/8-1:0];
            assign m_axis_fifo_12_tdata = dwconv_tdata[12][C_OUTPUT_FIFO_12_DMWIDTH-1:0];
            assign ap_fifo_oarg_12_full_n = full[12];
            assign write[12] = ap_fifo_oarg_12_write;
            assign din[12][C_OUTPUT_FIFO_12_WIDTH-1:0] = ap_fifo_oarg_12_din;
            assign tkeep[12] = {C_OUTPUT_FIFO_12_WIDTH/8{1'b1}};
            assign tstrb[12] = {C_OUTPUT_FIFO_12_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 13) begin
            assign dwconv_tready[13] = m_axis_fifo_13_tready;
            assign m_axis_fifo_13_tlast = dwconv_tlast[13];
            assign m_axis_fifo_13_tvalid = dwconv_tvalid[13];
            assign m_axis_fifo_13_tkeep = dwconv_tkeep[13][C_OUTPUT_FIFO_13_DMWIDTH/8-1:0];
            assign m_axis_fifo_13_tstrb = dwconv_tstrb[13][C_OUTPUT_FIFO_13_DMWIDTH/8-1:0];
            assign m_axis_fifo_13_tdata = dwconv_tdata[13][C_OUTPUT_FIFO_13_DMWIDTH-1:0];
            assign ap_fifo_oarg_13_full_n = full[13];
            assign write[13] = ap_fifo_oarg_13_write;
            assign din[13][C_OUTPUT_FIFO_13_WIDTH-1:0] = ap_fifo_oarg_13_din;
            assign tkeep[13] = {C_OUTPUT_FIFO_13_WIDTH/8{1'b1}};
            assign tstrb[13] = {C_OUTPUT_FIFO_13_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 14) begin
            assign dwconv_tready[14] = m_axis_fifo_14_tready;
            assign m_axis_fifo_14_tlast = dwconv_tlast[14];
            assign m_axis_fifo_14_tvalid = dwconv_tvalid[14];
            assign m_axis_fifo_14_tkeep = dwconv_tkeep[14][C_OUTPUT_FIFO_14_DMWIDTH/8-1:0];
            assign m_axis_fifo_14_tstrb = dwconv_tstrb[14][C_OUTPUT_FIFO_14_DMWIDTH/8-1:0];
            assign m_axis_fifo_14_tdata = dwconv_tdata[14][C_OUTPUT_FIFO_14_DMWIDTH-1:0];
            assign ap_fifo_oarg_14_full_n = full[14];
            assign write[14] = ap_fifo_oarg_14_write;
            assign din[14][C_OUTPUT_FIFO_14_WIDTH-1:0] = ap_fifo_oarg_14_din;
            assign tkeep[14] = {C_OUTPUT_FIFO_14_WIDTH/8{1'b1}};
            assign tstrb[14] = {C_OUTPUT_FIFO_14_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 15) begin
            assign dwconv_tready[15] = m_axis_fifo_15_tready;
            assign m_axis_fifo_15_tlast = dwconv_tlast[15];
            assign m_axis_fifo_15_tvalid = dwconv_tvalid[15];
            assign m_axis_fifo_15_tkeep = dwconv_tkeep[15][C_OUTPUT_FIFO_15_DMWIDTH/8-1:0];
            assign m_axis_fifo_15_tstrb = dwconv_tstrb[15][C_OUTPUT_FIFO_15_DMWIDTH/8-1:0];
            assign m_axis_fifo_15_tdata = dwconv_tdata[15][C_OUTPUT_FIFO_15_DMWIDTH-1:0];
            assign ap_fifo_oarg_15_full_n = full[15];
            assign write[15] = ap_fifo_oarg_15_write;
            assign din[15][C_OUTPUT_FIFO_15_WIDTH-1:0] = ap_fifo_oarg_15_din;
            assign tkeep[15] = {C_OUTPUT_FIFO_15_WIDTH/8{1'b1}};
            assign tstrb[15] = {C_OUTPUT_FIFO_15_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 16) begin
            assign dwconv_tready[16] = m_axis_fifo_16_tready;
            assign m_axis_fifo_16_tlast = dwconv_tlast[16];
            assign m_axis_fifo_16_tvalid = dwconv_tvalid[16];
            assign m_axis_fifo_16_tkeep = dwconv_tkeep[16][C_OUTPUT_FIFO_16_DMWIDTH/8-1:0];
            assign m_axis_fifo_16_tstrb = dwconv_tstrb[16][C_OUTPUT_FIFO_16_DMWIDTH/8-1:0];
            assign m_axis_fifo_16_tdata = dwconv_tdata[16][C_OUTPUT_FIFO_16_DMWIDTH-1:0];
            assign ap_fifo_oarg_16_full_n = full[16];
            assign write[16] = ap_fifo_oarg_16_write;
            assign din[16][C_OUTPUT_FIFO_16_WIDTH-1:0] = ap_fifo_oarg_16_din;
            assign tkeep[16] = {C_OUTPUT_FIFO_16_WIDTH/8{1'b1}};
            assign tstrb[16] = {C_OUTPUT_FIFO_16_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 17) begin
            assign dwconv_tready[17] = m_axis_fifo_17_tready;
            assign m_axis_fifo_17_tlast = dwconv_tlast[17];
            assign m_axis_fifo_17_tvalid = dwconv_tvalid[17];
            assign m_axis_fifo_17_tkeep = dwconv_tkeep[17][C_OUTPUT_FIFO_17_DMWIDTH/8-1:0];
            assign m_axis_fifo_17_tstrb = dwconv_tstrb[17][C_OUTPUT_FIFO_17_DMWIDTH/8-1:0];
            assign m_axis_fifo_17_tdata = dwconv_tdata[17][C_OUTPUT_FIFO_17_DMWIDTH-1:0];
            assign ap_fifo_oarg_17_full_n = full[17];
            assign write[17] = ap_fifo_oarg_17_write;
            assign din[17][C_OUTPUT_FIFO_17_WIDTH-1:0] = ap_fifo_oarg_17_din;
            assign tkeep[17] = {C_OUTPUT_FIFO_17_WIDTH/8{1'b1}};
            assign tstrb[17] = {C_OUTPUT_FIFO_17_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 18) begin
            assign dwconv_tready[18] = m_axis_fifo_18_tready;
            assign m_axis_fifo_18_tlast = dwconv_tlast[18];
            assign m_axis_fifo_18_tvalid = dwconv_tvalid[18];
            assign m_axis_fifo_18_tkeep = dwconv_tkeep[18][C_OUTPUT_FIFO_18_DMWIDTH/8-1:0];
            assign m_axis_fifo_18_tstrb = dwconv_tstrb[18][C_OUTPUT_FIFO_18_DMWIDTH/8-1:0];
            assign m_axis_fifo_18_tdata = dwconv_tdata[18][C_OUTPUT_FIFO_18_DMWIDTH-1:0];
            assign ap_fifo_oarg_18_full_n = full[18];
            assign write[18] = ap_fifo_oarg_18_write;
            assign din[18][C_OUTPUT_FIFO_18_WIDTH-1:0] = ap_fifo_oarg_18_din;
            assign tkeep[18] = {C_OUTPUT_FIFO_18_WIDTH/8{1'b1}};
            assign tstrb[18] = {C_OUTPUT_FIFO_18_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 19) begin
            assign dwconv_tready[19] = m_axis_fifo_19_tready;
            assign m_axis_fifo_19_tlast = dwconv_tlast[19];
            assign m_axis_fifo_19_tvalid = dwconv_tvalid[19];
            assign m_axis_fifo_19_tkeep = dwconv_tkeep[19][C_OUTPUT_FIFO_19_DMWIDTH/8-1:0];
            assign m_axis_fifo_19_tstrb = dwconv_tstrb[19][C_OUTPUT_FIFO_19_DMWIDTH/8-1:0];
            assign m_axis_fifo_19_tdata = dwconv_tdata[19][C_OUTPUT_FIFO_19_DMWIDTH-1:0];
            assign ap_fifo_oarg_19_full_n = full[19];
            assign write[19] = ap_fifo_oarg_19_write;
            assign din[19][C_OUTPUT_FIFO_19_WIDTH-1:0] = ap_fifo_oarg_19_din;
            assign tkeep[19] = {C_OUTPUT_FIFO_19_WIDTH/8{1'b1}};
            assign tstrb[19] = {C_OUTPUT_FIFO_19_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 20) begin
            assign dwconv_tready[20] = m_axis_fifo_20_tready;
            assign m_axis_fifo_20_tlast = dwconv_tlast[20];
            assign m_axis_fifo_20_tvalid = dwconv_tvalid[20];
            assign m_axis_fifo_20_tkeep = dwconv_tkeep[20][C_OUTPUT_FIFO_20_DMWIDTH/8-1:0];
            assign m_axis_fifo_20_tstrb = dwconv_tstrb[20][C_OUTPUT_FIFO_20_DMWIDTH/8-1:0];
            assign m_axis_fifo_20_tdata = dwconv_tdata[20][C_OUTPUT_FIFO_20_DMWIDTH-1:0];
            assign ap_fifo_oarg_20_full_n = full[20];
            assign write[20] = ap_fifo_oarg_20_write;
            assign din[20][C_OUTPUT_FIFO_20_WIDTH-1:0] = ap_fifo_oarg_20_din;
            assign tkeep[20] = {C_OUTPUT_FIFO_20_WIDTH/8{1'b1}};
            assign tstrb[20] = {C_OUTPUT_FIFO_20_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 21) begin
            assign dwconv_tready[21] = m_axis_fifo_21_tready;
            assign m_axis_fifo_21_tlast = dwconv_tlast[21];
            assign m_axis_fifo_21_tvalid = dwconv_tvalid[21];
            assign m_axis_fifo_21_tkeep = dwconv_tkeep[21][C_OUTPUT_FIFO_21_DMWIDTH/8-1:0];
            assign m_axis_fifo_21_tstrb = dwconv_tstrb[21][C_OUTPUT_FIFO_21_DMWIDTH/8-1:0];
            assign m_axis_fifo_21_tdata = dwconv_tdata[21][C_OUTPUT_FIFO_21_DMWIDTH-1:0];
            assign ap_fifo_oarg_21_full_n = full[21];
            assign write[21] = ap_fifo_oarg_21_write;
            assign din[21][C_OUTPUT_FIFO_21_WIDTH-1:0] = ap_fifo_oarg_21_din;
            assign tkeep[21] = {C_OUTPUT_FIFO_21_WIDTH/8{1'b1}};
            assign tstrb[21] = {C_OUTPUT_FIFO_21_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 22) begin
            assign dwconv_tready[22] = m_axis_fifo_22_tready;
            assign m_axis_fifo_22_tlast = dwconv_tlast[22];
            assign m_axis_fifo_22_tvalid = dwconv_tvalid[22];
            assign m_axis_fifo_22_tkeep = dwconv_tkeep[22][C_OUTPUT_FIFO_22_DMWIDTH/8-1:0];
            assign m_axis_fifo_22_tstrb = dwconv_tstrb[22][C_OUTPUT_FIFO_22_DMWIDTH/8-1:0];
            assign m_axis_fifo_22_tdata = dwconv_tdata[22][C_OUTPUT_FIFO_22_DMWIDTH-1:0];
            assign ap_fifo_oarg_22_full_n = full[22];
            assign write[22] = ap_fifo_oarg_22_write;
            assign din[22][C_OUTPUT_FIFO_22_WIDTH-1:0] = ap_fifo_oarg_22_din;
            assign tkeep[22] = {C_OUTPUT_FIFO_22_WIDTH/8{1'b1}};
            assign tstrb[22] = {C_OUTPUT_FIFO_22_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 23) begin
            assign dwconv_tready[23] = m_axis_fifo_23_tready;
            assign m_axis_fifo_23_tlast = dwconv_tlast[23];
            assign m_axis_fifo_23_tvalid = dwconv_tvalid[23];
            assign m_axis_fifo_23_tkeep = dwconv_tkeep[23][C_OUTPUT_FIFO_23_DMWIDTH/8-1:0];
            assign m_axis_fifo_23_tstrb = dwconv_tstrb[23][C_OUTPUT_FIFO_23_DMWIDTH/8-1:0];
            assign m_axis_fifo_23_tdata = dwconv_tdata[23][C_OUTPUT_FIFO_23_DMWIDTH-1:0];
            assign ap_fifo_oarg_23_full_n = full[23];
            assign write[23] = ap_fifo_oarg_23_write;
            assign din[23][C_OUTPUT_FIFO_23_WIDTH-1:0] = ap_fifo_oarg_23_din;
            assign tkeep[23] = {C_OUTPUT_FIFO_23_WIDTH/8{1'b1}};
            assign tstrb[23] = {C_OUTPUT_FIFO_23_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 24) begin
            assign dwconv_tready[24] = m_axis_fifo_24_tready;
            assign m_axis_fifo_24_tlast = dwconv_tlast[24];
            assign m_axis_fifo_24_tvalid = dwconv_tvalid[24];
            assign m_axis_fifo_24_tkeep = dwconv_tkeep[24][C_OUTPUT_FIFO_24_DMWIDTH/8-1:0];
            assign m_axis_fifo_24_tstrb = dwconv_tstrb[24][C_OUTPUT_FIFO_24_DMWIDTH/8-1:0];
            assign m_axis_fifo_24_tdata = dwconv_tdata[24][C_OUTPUT_FIFO_24_DMWIDTH-1:0];
            assign ap_fifo_oarg_24_full_n = full[24];
            assign write[24] = ap_fifo_oarg_24_write;
            assign din[24][C_OUTPUT_FIFO_24_WIDTH-1:0] = ap_fifo_oarg_24_din;
            assign tkeep[24] = {C_OUTPUT_FIFO_24_WIDTH/8{1'b1}};
            assign tstrb[24] = {C_OUTPUT_FIFO_24_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 25) begin
            assign dwconv_tready[25] = m_axis_fifo_25_tready;
            assign m_axis_fifo_25_tlast = dwconv_tlast[25];
            assign m_axis_fifo_25_tvalid = dwconv_tvalid[25];
            assign m_axis_fifo_25_tkeep = dwconv_tkeep[25][C_OUTPUT_FIFO_25_DMWIDTH/8-1:0];
            assign m_axis_fifo_25_tstrb = dwconv_tstrb[25][C_OUTPUT_FIFO_25_DMWIDTH/8-1:0];
            assign m_axis_fifo_25_tdata = dwconv_tdata[25][C_OUTPUT_FIFO_25_DMWIDTH-1:0];
            assign ap_fifo_oarg_25_full_n = full[25];
            assign write[25] = ap_fifo_oarg_25_write;
            assign din[25][C_OUTPUT_FIFO_25_WIDTH-1:0] = ap_fifo_oarg_25_din;
            assign tkeep[25] = {C_OUTPUT_FIFO_25_WIDTH/8{1'b1}};
            assign tstrb[25] = {C_OUTPUT_FIFO_25_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 26) begin
            assign dwconv_tready[26] = m_axis_fifo_26_tready;
            assign m_axis_fifo_26_tlast = dwconv_tlast[26];
            assign m_axis_fifo_26_tvalid = dwconv_tvalid[26];
            assign m_axis_fifo_26_tkeep = dwconv_tkeep[26][C_OUTPUT_FIFO_26_DMWIDTH/8-1:0];
            assign m_axis_fifo_26_tstrb = dwconv_tstrb[26][C_OUTPUT_FIFO_26_DMWIDTH/8-1:0];
            assign m_axis_fifo_26_tdata = dwconv_tdata[26][C_OUTPUT_FIFO_26_DMWIDTH-1:0];
            assign ap_fifo_oarg_26_full_n = full[26];
            assign write[26] = ap_fifo_oarg_26_write;
            assign din[26][C_OUTPUT_FIFO_26_WIDTH-1:0] = ap_fifo_oarg_26_din;
            assign tkeep[26] = {C_OUTPUT_FIFO_26_WIDTH/8{1'b1}};
            assign tstrb[26] = {C_OUTPUT_FIFO_26_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 27) begin
            assign dwconv_tready[27] = m_axis_fifo_27_tready;
            assign m_axis_fifo_27_tlast = dwconv_tlast[27];
            assign m_axis_fifo_27_tvalid = dwconv_tvalid[27];
            assign m_axis_fifo_27_tkeep = dwconv_tkeep[27][C_OUTPUT_FIFO_27_DMWIDTH/8-1:0];
            assign m_axis_fifo_27_tstrb = dwconv_tstrb[27][C_OUTPUT_FIFO_27_DMWIDTH/8-1:0];
            assign m_axis_fifo_27_tdata = dwconv_tdata[27][C_OUTPUT_FIFO_27_DMWIDTH-1:0];
            assign ap_fifo_oarg_27_full_n = full[27];
            assign write[27] = ap_fifo_oarg_27_write;
            assign din[27][C_OUTPUT_FIFO_27_WIDTH-1:0] = ap_fifo_oarg_27_din;
            assign tkeep[27] = {C_OUTPUT_FIFO_27_WIDTH/8{1'b1}};
            assign tstrb[27] = {C_OUTPUT_FIFO_27_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 28) begin
            assign dwconv_tready[28] = m_axis_fifo_28_tready;
            assign m_axis_fifo_28_tlast = dwconv_tlast[28];
            assign m_axis_fifo_28_tvalid = dwconv_tvalid[28];
            assign m_axis_fifo_28_tkeep = dwconv_tkeep[28][C_OUTPUT_FIFO_28_DMWIDTH/8-1:0];
            assign m_axis_fifo_28_tstrb = dwconv_tstrb[28][C_OUTPUT_FIFO_28_DMWIDTH/8-1:0];
            assign m_axis_fifo_28_tdata = dwconv_tdata[28][C_OUTPUT_FIFO_28_DMWIDTH-1:0];
            assign ap_fifo_oarg_28_full_n = full[28];
            assign write[28] = ap_fifo_oarg_28_write;
            assign din[28][C_OUTPUT_FIFO_28_WIDTH-1:0] = ap_fifo_oarg_28_din;
            assign tkeep[28] = {C_OUTPUT_FIFO_28_WIDTH/8{1'b1}};
            assign tstrb[28] = {C_OUTPUT_FIFO_28_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 29) begin
            assign dwconv_tready[29] = m_axis_fifo_29_tready;
            assign m_axis_fifo_29_tlast = dwconv_tlast[29];
            assign m_axis_fifo_29_tvalid = dwconv_tvalid[29];
            assign m_axis_fifo_29_tkeep = dwconv_tkeep[29][C_OUTPUT_FIFO_29_DMWIDTH/8-1:0];
            assign m_axis_fifo_29_tstrb = dwconv_tstrb[29][C_OUTPUT_FIFO_29_DMWIDTH/8-1:0];
            assign m_axis_fifo_29_tdata = dwconv_tdata[29][C_OUTPUT_FIFO_29_DMWIDTH-1:0];
            assign ap_fifo_oarg_29_full_n = full[29];
            assign write[29] = ap_fifo_oarg_29_write;
            assign din[29][C_OUTPUT_FIFO_29_WIDTH-1:0] = ap_fifo_oarg_29_din;
            assign tkeep[29] = {C_OUTPUT_FIFO_29_WIDTH/8{1'b1}};
            assign tstrb[29] = {C_OUTPUT_FIFO_29_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 30) begin
            assign dwconv_tready[30] = m_axis_fifo_30_tready;
            assign m_axis_fifo_30_tlast = dwconv_tlast[30];
            assign m_axis_fifo_30_tvalid = dwconv_tvalid[30];
            assign m_axis_fifo_30_tkeep = dwconv_tkeep[30][C_OUTPUT_FIFO_30_DMWIDTH/8-1:0];
            assign m_axis_fifo_30_tstrb = dwconv_tstrb[30][C_OUTPUT_FIFO_30_DMWIDTH/8-1:0];
            assign m_axis_fifo_30_tdata = dwconv_tdata[30][C_OUTPUT_FIFO_30_DMWIDTH-1:0];
            assign ap_fifo_oarg_30_full_n = full[30];
            assign write[30] = ap_fifo_oarg_30_write;
            assign din[30][C_OUTPUT_FIFO_30_WIDTH-1:0] = ap_fifo_oarg_30_din;
            assign tkeep[30] = {C_OUTPUT_FIFO_30_WIDTH/8{1'b1}};
            assign tstrb[30] = {C_OUTPUT_FIFO_30_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 31) begin
            assign dwconv_tready[31] = m_axis_fifo_31_tready;
            assign m_axis_fifo_31_tlast = dwconv_tlast[31];
            assign m_axis_fifo_31_tvalid = dwconv_tvalid[31];
            assign m_axis_fifo_31_tkeep = dwconv_tkeep[31][C_OUTPUT_FIFO_31_DMWIDTH/8-1:0];
            assign m_axis_fifo_31_tstrb = dwconv_tstrb[31][C_OUTPUT_FIFO_31_DMWIDTH/8-1:0];
            assign m_axis_fifo_31_tdata = dwconv_tdata[31][C_OUTPUT_FIFO_31_DMWIDTH-1:0];
            assign ap_fifo_oarg_31_full_n = full[31];
            assign write[31] = ap_fifo_oarg_31_write;
            assign din[31][C_OUTPUT_FIFO_31_WIDTH-1:0] = ap_fifo_oarg_31_din;
            assign tkeep[31] = {C_OUTPUT_FIFO_31_WIDTH/8{1'b1}};
            assign tstrb[31] = {C_OUTPUT_FIFO_31_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 32) begin
            assign dwconv_tready[32] = m_axis_fifo_32_tready;
            assign m_axis_fifo_32_tlast = dwconv_tlast[32];
            assign m_axis_fifo_32_tvalid = dwconv_tvalid[32];
            assign m_axis_fifo_32_tkeep = dwconv_tkeep[32][C_OUTPUT_FIFO_32_DMWIDTH/8-1:0];
            assign m_axis_fifo_32_tstrb = dwconv_tstrb[32][C_OUTPUT_FIFO_32_DMWIDTH/8-1:0];
            assign m_axis_fifo_32_tdata = dwconv_tdata[32][C_OUTPUT_FIFO_32_DMWIDTH-1:0];
            assign ap_fifo_oarg_32_full_n = full[32];
            assign write[32] = ap_fifo_oarg_32_write;
            assign din[32][C_OUTPUT_FIFO_32_WIDTH-1:0] = ap_fifo_oarg_32_din;
            assign tkeep[32] = {C_OUTPUT_FIFO_32_WIDTH/8{1'b1}};
            assign tstrb[32] = {C_OUTPUT_FIFO_32_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 33) begin
            assign dwconv_tready[33] = m_axis_fifo_33_tready;
            assign m_axis_fifo_33_tlast = dwconv_tlast[33];
            assign m_axis_fifo_33_tvalid = dwconv_tvalid[33];
            assign m_axis_fifo_33_tkeep = dwconv_tkeep[33][C_OUTPUT_FIFO_33_DMWIDTH/8-1:0];
            assign m_axis_fifo_33_tstrb = dwconv_tstrb[33][C_OUTPUT_FIFO_33_DMWIDTH/8-1:0];
            assign m_axis_fifo_33_tdata = dwconv_tdata[33][C_OUTPUT_FIFO_33_DMWIDTH-1:0];
            assign ap_fifo_oarg_33_full_n = full[33];
            assign write[33] = ap_fifo_oarg_33_write;
            assign din[33][C_OUTPUT_FIFO_33_WIDTH-1:0] = ap_fifo_oarg_33_din;
            assign tkeep[33] = {C_OUTPUT_FIFO_33_WIDTH/8{1'b1}};
            assign tstrb[33] = {C_OUTPUT_FIFO_33_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 34) begin
            assign dwconv_tready[34] = m_axis_fifo_34_tready;
            assign m_axis_fifo_34_tlast = dwconv_tlast[34];
            assign m_axis_fifo_34_tvalid = dwconv_tvalid[34];
            assign m_axis_fifo_34_tkeep = dwconv_tkeep[34][C_OUTPUT_FIFO_34_DMWIDTH/8-1:0];
            assign m_axis_fifo_34_tstrb = dwconv_tstrb[34][C_OUTPUT_FIFO_34_DMWIDTH/8-1:0];
            assign m_axis_fifo_34_tdata = dwconv_tdata[34][C_OUTPUT_FIFO_34_DMWIDTH-1:0];
            assign ap_fifo_oarg_34_full_n = full[34];
            assign write[34] = ap_fifo_oarg_34_write;
            assign din[34][C_OUTPUT_FIFO_34_WIDTH-1:0] = ap_fifo_oarg_34_din;
            assign tkeep[34] = {C_OUTPUT_FIFO_34_WIDTH/8{1'b1}};
            assign tstrb[34] = {C_OUTPUT_FIFO_34_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 35) begin
            assign dwconv_tready[35] = m_axis_fifo_35_tready;
            assign m_axis_fifo_35_tlast = dwconv_tlast[35];
            assign m_axis_fifo_35_tvalid = dwconv_tvalid[35];
            assign m_axis_fifo_35_tkeep = dwconv_tkeep[35][C_OUTPUT_FIFO_35_DMWIDTH/8-1:0];
            assign m_axis_fifo_35_tstrb = dwconv_tstrb[35][C_OUTPUT_FIFO_35_DMWIDTH/8-1:0];
            assign m_axis_fifo_35_tdata = dwconv_tdata[35][C_OUTPUT_FIFO_35_DMWIDTH-1:0];
            assign ap_fifo_oarg_35_full_n = full[35];
            assign write[35] = ap_fifo_oarg_35_write;
            assign din[35][C_OUTPUT_FIFO_35_WIDTH-1:0] = ap_fifo_oarg_35_din;
            assign tkeep[35] = {C_OUTPUT_FIFO_35_WIDTH/8{1'b1}};
            assign tstrb[35] = {C_OUTPUT_FIFO_35_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 36) begin
            assign dwconv_tready[36] = m_axis_fifo_36_tready;
            assign m_axis_fifo_36_tlast = dwconv_tlast[36];
            assign m_axis_fifo_36_tvalid = dwconv_tvalid[36];
            assign m_axis_fifo_36_tkeep = dwconv_tkeep[36][C_OUTPUT_FIFO_36_DMWIDTH/8-1:0];
            assign m_axis_fifo_36_tstrb = dwconv_tstrb[36][C_OUTPUT_FIFO_36_DMWIDTH/8-1:0];
            assign m_axis_fifo_36_tdata = dwconv_tdata[36][C_OUTPUT_FIFO_36_DMWIDTH-1:0];
            assign ap_fifo_oarg_36_full_n = full[36];
            assign write[36] = ap_fifo_oarg_36_write;
            assign din[36][C_OUTPUT_FIFO_36_WIDTH-1:0] = ap_fifo_oarg_36_din;
            assign tkeep[36] = {C_OUTPUT_FIFO_36_WIDTH/8{1'b1}};
            assign tstrb[36] = {C_OUTPUT_FIFO_36_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 37) begin
            assign dwconv_tready[37] = m_axis_fifo_37_tready;
            assign m_axis_fifo_37_tlast = dwconv_tlast[37];
            assign m_axis_fifo_37_tvalid = dwconv_tvalid[37];
            assign m_axis_fifo_37_tkeep = dwconv_tkeep[37][C_OUTPUT_FIFO_37_DMWIDTH/8-1:0];
            assign m_axis_fifo_37_tstrb = dwconv_tstrb[37][C_OUTPUT_FIFO_37_DMWIDTH/8-1:0];
            assign m_axis_fifo_37_tdata = dwconv_tdata[37][C_OUTPUT_FIFO_37_DMWIDTH-1:0];
            assign ap_fifo_oarg_37_full_n = full[37];
            assign write[37] = ap_fifo_oarg_37_write;
            assign din[37][C_OUTPUT_FIFO_37_WIDTH-1:0] = ap_fifo_oarg_37_din;
            assign tkeep[37] = {C_OUTPUT_FIFO_37_WIDTH/8{1'b1}};
            assign tstrb[37] = {C_OUTPUT_FIFO_37_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 38) begin
            assign dwconv_tready[38] = m_axis_fifo_38_tready;
            assign m_axis_fifo_38_tlast = dwconv_tlast[38];
            assign m_axis_fifo_38_tvalid = dwconv_tvalid[38];
            assign m_axis_fifo_38_tkeep = dwconv_tkeep[38][C_OUTPUT_FIFO_38_DMWIDTH/8-1:0];
            assign m_axis_fifo_38_tstrb = dwconv_tstrb[38][C_OUTPUT_FIFO_38_DMWIDTH/8-1:0];
            assign m_axis_fifo_38_tdata = dwconv_tdata[38][C_OUTPUT_FIFO_38_DMWIDTH-1:0];
            assign ap_fifo_oarg_38_full_n = full[38];
            assign write[38] = ap_fifo_oarg_38_write;
            assign din[38][C_OUTPUT_FIFO_38_WIDTH-1:0] = ap_fifo_oarg_38_din;
            assign tkeep[38] = {C_OUTPUT_FIFO_38_WIDTH/8{1'b1}};
            assign tstrb[38] = {C_OUTPUT_FIFO_38_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 39) begin
            assign dwconv_tready[39] = m_axis_fifo_39_tready;
            assign m_axis_fifo_39_tlast = dwconv_tlast[39];
            assign m_axis_fifo_39_tvalid = dwconv_tvalid[39];
            assign m_axis_fifo_39_tkeep = dwconv_tkeep[39][C_OUTPUT_FIFO_39_DMWIDTH/8-1:0];
            assign m_axis_fifo_39_tstrb = dwconv_tstrb[39][C_OUTPUT_FIFO_39_DMWIDTH/8-1:0];
            assign m_axis_fifo_39_tdata = dwconv_tdata[39][C_OUTPUT_FIFO_39_DMWIDTH-1:0];
            assign ap_fifo_oarg_39_full_n = full[39];
            assign write[39] = ap_fifo_oarg_39_write;
            assign din[39][C_OUTPUT_FIFO_39_WIDTH-1:0] = ap_fifo_oarg_39_din;
            assign tkeep[39] = {C_OUTPUT_FIFO_39_WIDTH/8{1'b1}};
            assign tstrb[39] = {C_OUTPUT_FIFO_39_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 40) begin
            assign dwconv_tready[40] = m_axis_fifo_40_tready;
            assign m_axis_fifo_40_tlast = dwconv_tlast[40];
            assign m_axis_fifo_40_tvalid = dwconv_tvalid[40];
            assign m_axis_fifo_40_tkeep = dwconv_tkeep[40][C_OUTPUT_FIFO_40_DMWIDTH/8-1:0];
            assign m_axis_fifo_40_tstrb = dwconv_tstrb[40][C_OUTPUT_FIFO_40_DMWIDTH/8-1:0];
            assign m_axis_fifo_40_tdata = dwconv_tdata[40][C_OUTPUT_FIFO_40_DMWIDTH-1:0];
            assign ap_fifo_oarg_40_full_n = full[40];
            assign write[40] = ap_fifo_oarg_40_write;
            assign din[40][C_OUTPUT_FIFO_40_WIDTH-1:0] = ap_fifo_oarg_40_din;
            assign tkeep[40] = {C_OUTPUT_FIFO_40_WIDTH/8{1'b1}};
            assign tstrb[40] = {C_OUTPUT_FIFO_40_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 41) begin
            assign dwconv_tready[41] = m_axis_fifo_41_tready;
            assign m_axis_fifo_41_tlast = dwconv_tlast[41];
            assign m_axis_fifo_41_tvalid = dwconv_tvalid[41];
            assign m_axis_fifo_41_tkeep = dwconv_tkeep[41][C_OUTPUT_FIFO_41_DMWIDTH/8-1:0];
            assign m_axis_fifo_41_tstrb = dwconv_tstrb[41][C_OUTPUT_FIFO_41_DMWIDTH/8-1:0];
            assign m_axis_fifo_41_tdata = dwconv_tdata[41][C_OUTPUT_FIFO_41_DMWIDTH-1:0];
            assign ap_fifo_oarg_41_full_n = full[41];
            assign write[41] = ap_fifo_oarg_41_write;
            assign din[41][C_OUTPUT_FIFO_41_WIDTH-1:0] = ap_fifo_oarg_41_din;
            assign tkeep[41] = {C_OUTPUT_FIFO_41_WIDTH/8{1'b1}};
            assign tstrb[41] = {C_OUTPUT_FIFO_41_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 42) begin
            assign dwconv_tready[42] = m_axis_fifo_42_tready;
            assign m_axis_fifo_42_tlast = dwconv_tlast[42];
            assign m_axis_fifo_42_tvalid = dwconv_tvalid[42];
            assign m_axis_fifo_42_tkeep = dwconv_tkeep[42][C_OUTPUT_FIFO_42_DMWIDTH/8-1:0];
            assign m_axis_fifo_42_tstrb = dwconv_tstrb[42][C_OUTPUT_FIFO_42_DMWIDTH/8-1:0];
            assign m_axis_fifo_42_tdata = dwconv_tdata[42][C_OUTPUT_FIFO_42_DMWIDTH-1:0];
            assign ap_fifo_oarg_42_full_n = full[42];
            assign write[42] = ap_fifo_oarg_42_write;
            assign din[42][C_OUTPUT_FIFO_42_WIDTH-1:0] = ap_fifo_oarg_42_din;
            assign tkeep[42] = {C_OUTPUT_FIFO_42_WIDTH/8{1'b1}};
            assign tstrb[42] = {C_OUTPUT_FIFO_42_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 43) begin
            assign dwconv_tready[43] = m_axis_fifo_43_tready;
            assign m_axis_fifo_43_tlast = dwconv_tlast[43];
            assign m_axis_fifo_43_tvalid = dwconv_tvalid[43];
            assign m_axis_fifo_43_tkeep = dwconv_tkeep[43][C_OUTPUT_FIFO_43_DMWIDTH/8-1:0];
            assign m_axis_fifo_43_tstrb = dwconv_tstrb[43][C_OUTPUT_FIFO_43_DMWIDTH/8-1:0];
            assign m_axis_fifo_43_tdata = dwconv_tdata[43][C_OUTPUT_FIFO_43_DMWIDTH-1:0];
            assign ap_fifo_oarg_43_full_n = full[43];
            assign write[43] = ap_fifo_oarg_43_write;
            assign din[43][C_OUTPUT_FIFO_43_WIDTH-1:0] = ap_fifo_oarg_43_din;
            assign tkeep[43] = {C_OUTPUT_FIFO_43_WIDTH/8{1'b1}};
            assign tstrb[43] = {C_OUTPUT_FIFO_43_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 44) begin
            assign dwconv_tready[44] = m_axis_fifo_44_tready;
            assign m_axis_fifo_44_tlast = dwconv_tlast[44];
            assign m_axis_fifo_44_tvalid = dwconv_tvalid[44];
            assign m_axis_fifo_44_tkeep = dwconv_tkeep[44][C_OUTPUT_FIFO_44_DMWIDTH/8-1:0];
            assign m_axis_fifo_44_tstrb = dwconv_tstrb[44][C_OUTPUT_FIFO_44_DMWIDTH/8-1:0];
            assign m_axis_fifo_44_tdata = dwconv_tdata[44][C_OUTPUT_FIFO_44_DMWIDTH-1:0];
            assign ap_fifo_oarg_44_full_n = full[44];
            assign write[44] = ap_fifo_oarg_44_write;
            assign din[44][C_OUTPUT_FIFO_44_WIDTH-1:0] = ap_fifo_oarg_44_din;
            assign tkeep[44] = {C_OUTPUT_FIFO_44_WIDTH/8{1'b1}};
            assign tstrb[44] = {C_OUTPUT_FIFO_44_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 45) begin
            assign dwconv_tready[45] = m_axis_fifo_45_tready;
            assign m_axis_fifo_45_tlast = dwconv_tlast[45];
            assign m_axis_fifo_45_tvalid = dwconv_tvalid[45];
            assign m_axis_fifo_45_tkeep = dwconv_tkeep[45][C_OUTPUT_FIFO_45_DMWIDTH/8-1:0];
            assign m_axis_fifo_45_tstrb = dwconv_tstrb[45][C_OUTPUT_FIFO_45_DMWIDTH/8-1:0];
            assign m_axis_fifo_45_tdata = dwconv_tdata[45][C_OUTPUT_FIFO_45_DMWIDTH-1:0];
            assign ap_fifo_oarg_45_full_n = full[45];
            assign write[45] = ap_fifo_oarg_45_write;
            assign din[45][C_OUTPUT_FIFO_45_WIDTH-1:0] = ap_fifo_oarg_45_din;
            assign tkeep[45] = {C_OUTPUT_FIFO_45_WIDTH/8{1'b1}};
            assign tstrb[45] = {C_OUTPUT_FIFO_45_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 46) begin
            assign dwconv_tready[46] = m_axis_fifo_46_tready;
            assign m_axis_fifo_46_tlast = dwconv_tlast[46];
            assign m_axis_fifo_46_tvalid = dwconv_tvalid[46];
            assign m_axis_fifo_46_tkeep = dwconv_tkeep[46][C_OUTPUT_FIFO_46_DMWIDTH/8-1:0];
            assign m_axis_fifo_46_tstrb = dwconv_tstrb[46][C_OUTPUT_FIFO_46_DMWIDTH/8-1:0];
            assign m_axis_fifo_46_tdata = dwconv_tdata[46][C_OUTPUT_FIFO_46_DMWIDTH-1:0];
            assign ap_fifo_oarg_46_full_n = full[46];
            assign write[46] = ap_fifo_oarg_46_write;
            assign din[46][C_OUTPUT_FIFO_46_WIDTH-1:0] = ap_fifo_oarg_46_din;
            assign tkeep[46] = {C_OUTPUT_FIFO_46_WIDTH/8{1'b1}};
            assign tstrb[46] = {C_OUTPUT_FIFO_46_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 47) begin
            assign dwconv_tready[47] = m_axis_fifo_47_tready;
            assign m_axis_fifo_47_tlast = dwconv_tlast[47];
            assign m_axis_fifo_47_tvalid = dwconv_tvalid[47];
            assign m_axis_fifo_47_tkeep = dwconv_tkeep[47][C_OUTPUT_FIFO_47_DMWIDTH/8-1:0];
            assign m_axis_fifo_47_tstrb = dwconv_tstrb[47][C_OUTPUT_FIFO_47_DMWIDTH/8-1:0];
            assign m_axis_fifo_47_tdata = dwconv_tdata[47][C_OUTPUT_FIFO_47_DMWIDTH-1:0];
            assign ap_fifo_oarg_47_full_n = full[47];
            assign write[47] = ap_fifo_oarg_47_write;
            assign din[47][C_OUTPUT_FIFO_47_WIDTH-1:0] = ap_fifo_oarg_47_din;
            assign tkeep[47] = {C_OUTPUT_FIFO_47_WIDTH/8{1'b1}};
            assign tstrb[47] = {C_OUTPUT_FIFO_47_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 48) begin
            assign dwconv_tready[48] = m_axis_fifo_48_tready;
            assign m_axis_fifo_48_tlast = dwconv_tlast[48];
            assign m_axis_fifo_48_tvalid = dwconv_tvalid[48];
            assign m_axis_fifo_48_tkeep = dwconv_tkeep[48][C_OUTPUT_FIFO_48_DMWIDTH/8-1:0];
            assign m_axis_fifo_48_tstrb = dwconv_tstrb[48][C_OUTPUT_FIFO_48_DMWIDTH/8-1:0];
            assign m_axis_fifo_48_tdata = dwconv_tdata[48][C_OUTPUT_FIFO_48_DMWIDTH-1:0];
            assign ap_fifo_oarg_48_full_n = full[48];
            assign write[48] = ap_fifo_oarg_48_write;
            assign din[48][C_OUTPUT_FIFO_48_WIDTH-1:0] = ap_fifo_oarg_48_din;
            assign tkeep[48] = {C_OUTPUT_FIFO_48_WIDTH/8{1'b1}};
            assign tstrb[48] = {C_OUTPUT_FIFO_48_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 49) begin
            assign dwconv_tready[49] = m_axis_fifo_49_tready;
            assign m_axis_fifo_49_tlast = dwconv_tlast[49];
            assign m_axis_fifo_49_tvalid = dwconv_tvalid[49];
            assign m_axis_fifo_49_tkeep = dwconv_tkeep[49][C_OUTPUT_FIFO_49_DMWIDTH/8-1:0];
            assign m_axis_fifo_49_tstrb = dwconv_tstrb[49][C_OUTPUT_FIFO_49_DMWIDTH/8-1:0];
            assign m_axis_fifo_49_tdata = dwconv_tdata[49][C_OUTPUT_FIFO_49_DMWIDTH-1:0];
            assign ap_fifo_oarg_49_full_n = full[49];
            assign write[49] = ap_fifo_oarg_49_write;
            assign din[49][C_OUTPUT_FIFO_49_WIDTH-1:0] = ap_fifo_oarg_49_din;
            assign tkeep[49] = {C_OUTPUT_FIFO_49_WIDTH/8{1'b1}};
            assign tstrb[49] = {C_OUTPUT_FIFO_49_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 50) begin
            assign dwconv_tready[50] = m_axis_fifo_50_tready;
            assign m_axis_fifo_50_tlast = dwconv_tlast[50];
            assign m_axis_fifo_50_tvalid = dwconv_tvalid[50];
            assign m_axis_fifo_50_tkeep = dwconv_tkeep[50][C_OUTPUT_FIFO_50_DMWIDTH/8-1:0];
            assign m_axis_fifo_50_tstrb = dwconv_tstrb[50][C_OUTPUT_FIFO_50_DMWIDTH/8-1:0];
            assign m_axis_fifo_50_tdata = dwconv_tdata[50][C_OUTPUT_FIFO_50_DMWIDTH-1:0];
            assign ap_fifo_oarg_50_full_n = full[50];
            assign write[50] = ap_fifo_oarg_50_write;
            assign din[50][C_OUTPUT_FIFO_50_WIDTH-1:0] = ap_fifo_oarg_50_din;
            assign tkeep[50] = {C_OUTPUT_FIFO_50_WIDTH/8{1'b1}};
            assign tstrb[50] = {C_OUTPUT_FIFO_50_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 51) begin
            assign dwconv_tready[51] = m_axis_fifo_51_tready;
            assign m_axis_fifo_51_tlast = dwconv_tlast[51];
            assign m_axis_fifo_51_tvalid = dwconv_tvalid[51];
            assign m_axis_fifo_51_tkeep = dwconv_tkeep[51][C_OUTPUT_FIFO_51_DMWIDTH/8-1:0];
            assign m_axis_fifo_51_tstrb = dwconv_tstrb[51][C_OUTPUT_FIFO_51_DMWIDTH/8-1:0];
            assign m_axis_fifo_51_tdata = dwconv_tdata[51][C_OUTPUT_FIFO_51_DMWIDTH-1:0];
            assign ap_fifo_oarg_51_full_n = full[51];
            assign write[51] = ap_fifo_oarg_51_write;
            assign din[51][C_OUTPUT_FIFO_51_WIDTH-1:0] = ap_fifo_oarg_51_din;
            assign tkeep[51] = {C_OUTPUT_FIFO_51_WIDTH/8{1'b1}};
            assign tstrb[51] = {C_OUTPUT_FIFO_51_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 52) begin
            assign dwconv_tready[52] = m_axis_fifo_52_tready;
            assign m_axis_fifo_52_tlast = dwconv_tlast[52];
            assign m_axis_fifo_52_tvalid = dwconv_tvalid[52];
            assign m_axis_fifo_52_tkeep = dwconv_tkeep[52][C_OUTPUT_FIFO_52_DMWIDTH/8-1:0];
            assign m_axis_fifo_52_tstrb = dwconv_tstrb[52][C_OUTPUT_FIFO_52_DMWIDTH/8-1:0];
            assign m_axis_fifo_52_tdata = dwconv_tdata[52][C_OUTPUT_FIFO_52_DMWIDTH-1:0];
            assign ap_fifo_oarg_52_full_n = full[52];
            assign write[52] = ap_fifo_oarg_52_write;
            assign din[52][C_OUTPUT_FIFO_52_WIDTH-1:0] = ap_fifo_oarg_52_din;
            assign tkeep[52] = {C_OUTPUT_FIFO_52_WIDTH/8{1'b1}};
            assign tstrb[52] = {C_OUTPUT_FIFO_52_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 53) begin
            assign dwconv_tready[53] = m_axis_fifo_53_tready;
            assign m_axis_fifo_53_tlast = dwconv_tlast[53];
            assign m_axis_fifo_53_tvalid = dwconv_tvalid[53];
            assign m_axis_fifo_53_tkeep = dwconv_tkeep[53][C_OUTPUT_FIFO_53_DMWIDTH/8-1:0];
            assign m_axis_fifo_53_tstrb = dwconv_tstrb[53][C_OUTPUT_FIFO_53_DMWIDTH/8-1:0];
            assign m_axis_fifo_53_tdata = dwconv_tdata[53][C_OUTPUT_FIFO_53_DMWIDTH-1:0];
            assign ap_fifo_oarg_53_full_n = full[53];
            assign write[53] = ap_fifo_oarg_53_write;
            assign din[53][C_OUTPUT_FIFO_53_WIDTH-1:0] = ap_fifo_oarg_53_din;
            assign tkeep[53] = {C_OUTPUT_FIFO_53_WIDTH/8{1'b1}};
            assign tstrb[53] = {C_OUTPUT_FIFO_53_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 54) begin
            assign dwconv_tready[54] = m_axis_fifo_54_tready;
            assign m_axis_fifo_54_tlast = dwconv_tlast[54];
            assign m_axis_fifo_54_tvalid = dwconv_tvalid[54];
            assign m_axis_fifo_54_tkeep = dwconv_tkeep[54][C_OUTPUT_FIFO_54_DMWIDTH/8-1:0];
            assign m_axis_fifo_54_tstrb = dwconv_tstrb[54][C_OUTPUT_FIFO_54_DMWIDTH/8-1:0];
            assign m_axis_fifo_54_tdata = dwconv_tdata[54][C_OUTPUT_FIFO_54_DMWIDTH-1:0];
            assign ap_fifo_oarg_54_full_n = full[54];
            assign write[54] = ap_fifo_oarg_54_write;
            assign din[54][C_OUTPUT_FIFO_54_WIDTH-1:0] = ap_fifo_oarg_54_din;
            assign tkeep[54] = {C_OUTPUT_FIFO_54_WIDTH/8{1'b1}};
            assign tstrb[54] = {C_OUTPUT_FIFO_54_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 55) begin
            assign dwconv_tready[55] = m_axis_fifo_55_tready;
            assign m_axis_fifo_55_tlast = dwconv_tlast[55];
            assign m_axis_fifo_55_tvalid = dwconv_tvalid[55];
            assign m_axis_fifo_55_tkeep = dwconv_tkeep[55][C_OUTPUT_FIFO_55_DMWIDTH/8-1:0];
            assign m_axis_fifo_55_tstrb = dwconv_tstrb[55][C_OUTPUT_FIFO_55_DMWIDTH/8-1:0];
            assign m_axis_fifo_55_tdata = dwconv_tdata[55][C_OUTPUT_FIFO_55_DMWIDTH-1:0];
            assign ap_fifo_oarg_55_full_n = full[55];
            assign write[55] = ap_fifo_oarg_55_write;
            assign din[55][C_OUTPUT_FIFO_55_WIDTH-1:0] = ap_fifo_oarg_55_din;
            assign tkeep[55] = {C_OUTPUT_FIFO_55_WIDTH/8{1'b1}};
            assign tstrb[55] = {C_OUTPUT_FIFO_55_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 56) begin
            assign dwconv_tready[56] = m_axis_fifo_56_tready;
            assign m_axis_fifo_56_tlast = dwconv_tlast[56];
            assign m_axis_fifo_56_tvalid = dwconv_tvalid[56];
            assign m_axis_fifo_56_tkeep = dwconv_tkeep[56][C_OUTPUT_FIFO_56_DMWIDTH/8-1:0];
            assign m_axis_fifo_56_tstrb = dwconv_tstrb[56][C_OUTPUT_FIFO_56_DMWIDTH/8-1:0];
            assign m_axis_fifo_56_tdata = dwconv_tdata[56][C_OUTPUT_FIFO_56_DMWIDTH-1:0];
            assign ap_fifo_oarg_56_full_n = full[56];
            assign write[56] = ap_fifo_oarg_56_write;
            assign din[56][C_OUTPUT_FIFO_56_WIDTH-1:0] = ap_fifo_oarg_56_din;
            assign tkeep[56] = {C_OUTPUT_FIFO_56_WIDTH/8{1'b1}};
            assign tstrb[56] = {C_OUTPUT_FIFO_56_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 57) begin
            assign dwconv_tready[57] = m_axis_fifo_57_tready;
            assign m_axis_fifo_57_tlast = dwconv_tlast[57];
            assign m_axis_fifo_57_tvalid = dwconv_tvalid[57];
            assign m_axis_fifo_57_tkeep = dwconv_tkeep[57][C_OUTPUT_FIFO_57_DMWIDTH/8-1:0];
            assign m_axis_fifo_57_tstrb = dwconv_tstrb[57][C_OUTPUT_FIFO_57_DMWIDTH/8-1:0];
            assign m_axis_fifo_57_tdata = dwconv_tdata[57][C_OUTPUT_FIFO_57_DMWIDTH-1:0];
            assign ap_fifo_oarg_57_full_n = full[57];
            assign write[57] = ap_fifo_oarg_57_write;
            assign din[57][C_OUTPUT_FIFO_57_WIDTH-1:0] = ap_fifo_oarg_57_din;
            assign tkeep[57] = {C_OUTPUT_FIFO_57_WIDTH/8{1'b1}};
            assign tstrb[57] = {C_OUTPUT_FIFO_57_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 58) begin
            assign dwconv_tready[58] = m_axis_fifo_58_tready;
            assign m_axis_fifo_58_tlast = dwconv_tlast[58];
            assign m_axis_fifo_58_tvalid = dwconv_tvalid[58];
            assign m_axis_fifo_58_tkeep = dwconv_tkeep[58][C_OUTPUT_FIFO_58_DMWIDTH/8-1:0];
            assign m_axis_fifo_58_tstrb = dwconv_tstrb[58][C_OUTPUT_FIFO_58_DMWIDTH/8-1:0];
            assign m_axis_fifo_58_tdata = dwconv_tdata[58][C_OUTPUT_FIFO_58_DMWIDTH-1:0];
            assign ap_fifo_oarg_58_full_n = full[58];
            assign write[58] = ap_fifo_oarg_58_write;
            assign din[58][C_OUTPUT_FIFO_58_WIDTH-1:0] = ap_fifo_oarg_58_din;
            assign tkeep[58] = {C_OUTPUT_FIFO_58_WIDTH/8{1'b1}};
            assign tstrb[58] = {C_OUTPUT_FIFO_58_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 59) begin
            assign dwconv_tready[59] = m_axis_fifo_59_tready;
            assign m_axis_fifo_59_tlast = dwconv_tlast[59];
            assign m_axis_fifo_59_tvalid = dwconv_tvalid[59];
            assign m_axis_fifo_59_tkeep = dwconv_tkeep[59][C_OUTPUT_FIFO_59_DMWIDTH/8-1:0];
            assign m_axis_fifo_59_tstrb = dwconv_tstrb[59][C_OUTPUT_FIFO_59_DMWIDTH/8-1:0];
            assign m_axis_fifo_59_tdata = dwconv_tdata[59][C_OUTPUT_FIFO_59_DMWIDTH-1:0];
            assign ap_fifo_oarg_59_full_n = full[59];
            assign write[59] = ap_fifo_oarg_59_write;
            assign din[59][C_OUTPUT_FIFO_59_WIDTH-1:0] = ap_fifo_oarg_59_din;
            assign tkeep[59] = {C_OUTPUT_FIFO_59_WIDTH/8{1'b1}};
            assign tstrb[59] = {C_OUTPUT_FIFO_59_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 60) begin
            assign dwconv_tready[60] = m_axis_fifo_60_tready;
            assign m_axis_fifo_60_tlast = dwconv_tlast[60];
            assign m_axis_fifo_60_tvalid = dwconv_tvalid[60];
            assign m_axis_fifo_60_tkeep = dwconv_tkeep[60][C_OUTPUT_FIFO_60_DMWIDTH/8-1:0];
            assign m_axis_fifo_60_tstrb = dwconv_tstrb[60][C_OUTPUT_FIFO_60_DMWIDTH/8-1:0];
            assign m_axis_fifo_60_tdata = dwconv_tdata[60][C_OUTPUT_FIFO_60_DMWIDTH-1:0];
            assign ap_fifo_oarg_60_full_n = full[60];
            assign write[60] = ap_fifo_oarg_60_write;
            assign din[60][C_OUTPUT_FIFO_60_WIDTH-1:0] = ap_fifo_oarg_60_din;
            assign tkeep[60] = {C_OUTPUT_FIFO_60_WIDTH/8{1'b1}};
            assign tstrb[60] = {C_OUTPUT_FIFO_60_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 61) begin
            assign dwconv_tready[61] = m_axis_fifo_61_tready;
            assign m_axis_fifo_61_tlast = dwconv_tlast[61];
            assign m_axis_fifo_61_tvalid = dwconv_tvalid[61];
            assign m_axis_fifo_61_tkeep = dwconv_tkeep[61][C_OUTPUT_FIFO_61_DMWIDTH/8-1:0];
            assign m_axis_fifo_61_tstrb = dwconv_tstrb[61][C_OUTPUT_FIFO_61_DMWIDTH/8-1:0];
            assign m_axis_fifo_61_tdata = dwconv_tdata[61][C_OUTPUT_FIFO_61_DMWIDTH-1:0];
            assign ap_fifo_oarg_61_full_n = full[61];
            assign write[61] = ap_fifo_oarg_61_write;
            assign din[61][C_OUTPUT_FIFO_61_WIDTH-1:0] = ap_fifo_oarg_61_din;
            assign tkeep[61] = {C_OUTPUT_FIFO_61_WIDTH/8{1'b1}};
            assign tstrb[61] = {C_OUTPUT_FIFO_61_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 62) begin
            assign dwconv_tready[62] = m_axis_fifo_62_tready;
            assign m_axis_fifo_62_tlast = dwconv_tlast[62];
            assign m_axis_fifo_62_tvalid = dwconv_tvalid[62];
            assign m_axis_fifo_62_tkeep = dwconv_tkeep[62][C_OUTPUT_FIFO_62_DMWIDTH/8-1:0];
            assign m_axis_fifo_62_tstrb = dwconv_tstrb[62][C_OUTPUT_FIFO_62_DMWIDTH/8-1:0];
            assign m_axis_fifo_62_tdata = dwconv_tdata[62][C_OUTPUT_FIFO_62_DMWIDTH-1:0];
            assign ap_fifo_oarg_62_full_n = full[62];
            assign write[62] = ap_fifo_oarg_62_write;
            assign din[62][C_OUTPUT_FIFO_62_WIDTH-1:0] = ap_fifo_oarg_62_din;
            assign tkeep[62] = {C_OUTPUT_FIFO_62_WIDTH/8{1'b1}};
            assign tstrb[62] = {C_OUTPUT_FIFO_62_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 63) begin
            assign dwconv_tready[63] = m_axis_fifo_63_tready;
            assign m_axis_fifo_63_tlast = dwconv_tlast[63];
            assign m_axis_fifo_63_tvalid = dwconv_tvalid[63];
            assign m_axis_fifo_63_tkeep = dwconv_tkeep[63][C_OUTPUT_FIFO_63_DMWIDTH/8-1:0];
            assign m_axis_fifo_63_tstrb = dwconv_tstrb[63][C_OUTPUT_FIFO_63_DMWIDTH/8-1:0];
            assign m_axis_fifo_63_tdata = dwconv_tdata[63][C_OUTPUT_FIFO_63_DMWIDTH-1:0];
            assign ap_fifo_oarg_63_full_n = full[63];
            assign write[63] = ap_fifo_oarg_63_write;
            assign din[63][C_OUTPUT_FIFO_63_WIDTH-1:0] = ap_fifo_oarg_63_din;
            assign tkeep[63] = {C_OUTPUT_FIFO_63_WIDTH/8{1'b1}};
            assign tstrb[63] = {C_OUTPUT_FIFO_63_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 64) begin
            assign dwconv_tready[64] = m_axis_fifo_64_tready;
            assign m_axis_fifo_64_tlast = dwconv_tlast[64];
            assign m_axis_fifo_64_tvalid = dwconv_tvalid[64];
            assign m_axis_fifo_64_tkeep = dwconv_tkeep[64][C_OUTPUT_FIFO_64_DMWIDTH/8-1:0];
            assign m_axis_fifo_64_tstrb = dwconv_tstrb[64][C_OUTPUT_FIFO_64_DMWIDTH/8-1:0];
            assign m_axis_fifo_64_tdata = dwconv_tdata[64][C_OUTPUT_FIFO_64_DMWIDTH-1:0];
            assign ap_fifo_oarg_64_full_n = full[64];
            assign write[64] = ap_fifo_oarg_64_write;
            assign din[64][C_OUTPUT_FIFO_64_WIDTH-1:0] = ap_fifo_oarg_64_din;
            assign tkeep[64] = {C_OUTPUT_FIFO_64_WIDTH/8{1'b1}};
            assign tstrb[64] = {C_OUTPUT_FIFO_64_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 65) begin
            assign dwconv_tready[65] = m_axis_fifo_65_tready;
            assign m_axis_fifo_65_tlast = dwconv_tlast[65];
            assign m_axis_fifo_65_tvalid = dwconv_tvalid[65];
            assign m_axis_fifo_65_tkeep = dwconv_tkeep[65][C_OUTPUT_FIFO_65_DMWIDTH/8-1:0];
            assign m_axis_fifo_65_tstrb = dwconv_tstrb[65][C_OUTPUT_FIFO_65_DMWIDTH/8-1:0];
            assign m_axis_fifo_65_tdata = dwconv_tdata[65][C_OUTPUT_FIFO_65_DMWIDTH-1:0];
            assign ap_fifo_oarg_65_full_n = full[65];
            assign write[65] = ap_fifo_oarg_65_write;
            assign din[65][C_OUTPUT_FIFO_65_WIDTH-1:0] = ap_fifo_oarg_65_din;
            assign tkeep[65] = {C_OUTPUT_FIFO_65_WIDTH/8{1'b1}};
            assign tstrb[65] = {C_OUTPUT_FIFO_65_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 66) begin
            assign dwconv_tready[66] = m_axis_fifo_66_tready;
            assign m_axis_fifo_66_tlast = dwconv_tlast[66];
            assign m_axis_fifo_66_tvalid = dwconv_tvalid[66];
            assign m_axis_fifo_66_tkeep = dwconv_tkeep[66][C_OUTPUT_FIFO_66_DMWIDTH/8-1:0];
            assign m_axis_fifo_66_tstrb = dwconv_tstrb[66][C_OUTPUT_FIFO_66_DMWIDTH/8-1:0];
            assign m_axis_fifo_66_tdata = dwconv_tdata[66][C_OUTPUT_FIFO_66_DMWIDTH-1:0];
            assign ap_fifo_oarg_66_full_n = full[66];
            assign write[66] = ap_fifo_oarg_66_write;
            assign din[66][C_OUTPUT_FIFO_66_WIDTH-1:0] = ap_fifo_oarg_66_din;
            assign tkeep[66] = {C_OUTPUT_FIFO_66_WIDTH/8{1'b1}};
            assign tstrb[66] = {C_OUTPUT_FIFO_66_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 67) begin
            assign dwconv_tready[67] = m_axis_fifo_67_tready;
            assign m_axis_fifo_67_tlast = dwconv_tlast[67];
            assign m_axis_fifo_67_tvalid = dwconv_tvalid[67];
            assign m_axis_fifo_67_tkeep = dwconv_tkeep[67][C_OUTPUT_FIFO_67_DMWIDTH/8-1:0];
            assign m_axis_fifo_67_tstrb = dwconv_tstrb[67][C_OUTPUT_FIFO_67_DMWIDTH/8-1:0];
            assign m_axis_fifo_67_tdata = dwconv_tdata[67][C_OUTPUT_FIFO_67_DMWIDTH-1:0];
            assign ap_fifo_oarg_67_full_n = full[67];
            assign write[67] = ap_fifo_oarg_67_write;
            assign din[67][C_OUTPUT_FIFO_67_WIDTH-1:0] = ap_fifo_oarg_67_din;
            assign tkeep[67] = {C_OUTPUT_FIFO_67_WIDTH/8{1'b1}};
            assign tstrb[67] = {C_OUTPUT_FIFO_67_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 68) begin
            assign dwconv_tready[68] = m_axis_fifo_68_tready;
            assign m_axis_fifo_68_tlast = dwconv_tlast[68];
            assign m_axis_fifo_68_tvalid = dwconv_tvalid[68];
            assign m_axis_fifo_68_tkeep = dwconv_tkeep[68][C_OUTPUT_FIFO_68_DMWIDTH/8-1:0];
            assign m_axis_fifo_68_tstrb = dwconv_tstrb[68][C_OUTPUT_FIFO_68_DMWIDTH/8-1:0];
            assign m_axis_fifo_68_tdata = dwconv_tdata[68][C_OUTPUT_FIFO_68_DMWIDTH-1:0];
            assign ap_fifo_oarg_68_full_n = full[68];
            assign write[68] = ap_fifo_oarg_68_write;
            assign din[68][C_OUTPUT_FIFO_68_WIDTH-1:0] = ap_fifo_oarg_68_din;
            assign tkeep[68] = {C_OUTPUT_FIFO_68_WIDTH/8{1'b1}};
            assign tstrb[68] = {C_OUTPUT_FIFO_68_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 69) begin
            assign dwconv_tready[69] = m_axis_fifo_69_tready;
            assign m_axis_fifo_69_tlast = dwconv_tlast[69];
            assign m_axis_fifo_69_tvalid = dwconv_tvalid[69];
            assign m_axis_fifo_69_tkeep = dwconv_tkeep[69][C_OUTPUT_FIFO_69_DMWIDTH/8-1:0];
            assign m_axis_fifo_69_tstrb = dwconv_tstrb[69][C_OUTPUT_FIFO_69_DMWIDTH/8-1:0];
            assign m_axis_fifo_69_tdata = dwconv_tdata[69][C_OUTPUT_FIFO_69_DMWIDTH-1:0];
            assign ap_fifo_oarg_69_full_n = full[69];
            assign write[69] = ap_fifo_oarg_69_write;
            assign din[69][C_OUTPUT_FIFO_69_WIDTH-1:0] = ap_fifo_oarg_69_din;
            assign tkeep[69] = {C_OUTPUT_FIFO_69_WIDTH/8{1'b1}};
            assign tstrb[69] = {C_OUTPUT_FIFO_69_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 70) begin
            assign dwconv_tready[70] = m_axis_fifo_70_tready;
            assign m_axis_fifo_70_tlast = dwconv_tlast[70];
            assign m_axis_fifo_70_tvalid = dwconv_tvalid[70];
            assign m_axis_fifo_70_tkeep = dwconv_tkeep[70][C_OUTPUT_FIFO_70_DMWIDTH/8-1:0];
            assign m_axis_fifo_70_tstrb = dwconv_tstrb[70][C_OUTPUT_FIFO_70_DMWIDTH/8-1:0];
            assign m_axis_fifo_70_tdata = dwconv_tdata[70][C_OUTPUT_FIFO_70_DMWIDTH-1:0];
            assign ap_fifo_oarg_70_full_n = full[70];
            assign write[70] = ap_fifo_oarg_70_write;
            assign din[70][C_OUTPUT_FIFO_70_WIDTH-1:0] = ap_fifo_oarg_70_din;
            assign tkeep[70] = {C_OUTPUT_FIFO_70_WIDTH/8{1'b1}};
            assign tstrb[70] = {C_OUTPUT_FIFO_70_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 71) begin
            assign dwconv_tready[71] = m_axis_fifo_71_tready;
            assign m_axis_fifo_71_tlast = dwconv_tlast[71];
            assign m_axis_fifo_71_tvalid = dwconv_tvalid[71];
            assign m_axis_fifo_71_tkeep = dwconv_tkeep[71][C_OUTPUT_FIFO_71_DMWIDTH/8-1:0];
            assign m_axis_fifo_71_tstrb = dwconv_tstrb[71][C_OUTPUT_FIFO_71_DMWIDTH/8-1:0];
            assign m_axis_fifo_71_tdata = dwconv_tdata[71][C_OUTPUT_FIFO_71_DMWIDTH-1:0];
            assign ap_fifo_oarg_71_full_n = full[71];
            assign write[71] = ap_fifo_oarg_71_write;
            assign din[71][C_OUTPUT_FIFO_71_WIDTH-1:0] = ap_fifo_oarg_71_din;
            assign tkeep[71] = {C_OUTPUT_FIFO_71_WIDTH/8{1'b1}};
            assign tstrb[71] = {C_OUTPUT_FIFO_71_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 72) begin
            assign dwconv_tready[72] = m_axis_fifo_72_tready;
            assign m_axis_fifo_72_tlast = dwconv_tlast[72];
            assign m_axis_fifo_72_tvalid = dwconv_tvalid[72];
            assign m_axis_fifo_72_tkeep = dwconv_tkeep[72][C_OUTPUT_FIFO_72_DMWIDTH/8-1:0];
            assign m_axis_fifo_72_tstrb = dwconv_tstrb[72][C_OUTPUT_FIFO_72_DMWIDTH/8-1:0];
            assign m_axis_fifo_72_tdata = dwconv_tdata[72][C_OUTPUT_FIFO_72_DMWIDTH-1:0];
            assign ap_fifo_oarg_72_full_n = full[72];
            assign write[72] = ap_fifo_oarg_72_write;
            assign din[72][C_OUTPUT_FIFO_72_WIDTH-1:0] = ap_fifo_oarg_72_din;
            assign tkeep[72] = {C_OUTPUT_FIFO_72_WIDTH/8{1'b1}};
            assign tstrb[72] = {C_OUTPUT_FIFO_72_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 73) begin
            assign dwconv_tready[73] = m_axis_fifo_73_tready;
            assign m_axis_fifo_73_tlast = dwconv_tlast[73];
            assign m_axis_fifo_73_tvalid = dwconv_tvalid[73];
            assign m_axis_fifo_73_tkeep = dwconv_tkeep[73][C_OUTPUT_FIFO_73_DMWIDTH/8-1:0];
            assign m_axis_fifo_73_tstrb = dwconv_tstrb[73][C_OUTPUT_FIFO_73_DMWIDTH/8-1:0];
            assign m_axis_fifo_73_tdata = dwconv_tdata[73][C_OUTPUT_FIFO_73_DMWIDTH-1:0];
            assign ap_fifo_oarg_73_full_n = full[73];
            assign write[73] = ap_fifo_oarg_73_write;
            assign din[73][C_OUTPUT_FIFO_73_WIDTH-1:0] = ap_fifo_oarg_73_din;
            assign tkeep[73] = {C_OUTPUT_FIFO_73_WIDTH/8{1'b1}};
            assign tstrb[73] = {C_OUTPUT_FIFO_73_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 74) begin
            assign dwconv_tready[74] = m_axis_fifo_74_tready;
            assign m_axis_fifo_74_tlast = dwconv_tlast[74];
            assign m_axis_fifo_74_tvalid = dwconv_tvalid[74];
            assign m_axis_fifo_74_tkeep = dwconv_tkeep[74][C_OUTPUT_FIFO_74_DMWIDTH/8-1:0];
            assign m_axis_fifo_74_tstrb = dwconv_tstrb[74][C_OUTPUT_FIFO_74_DMWIDTH/8-1:0];
            assign m_axis_fifo_74_tdata = dwconv_tdata[74][C_OUTPUT_FIFO_74_DMWIDTH-1:0];
            assign ap_fifo_oarg_74_full_n = full[74];
            assign write[74] = ap_fifo_oarg_74_write;
            assign din[74][C_OUTPUT_FIFO_74_WIDTH-1:0] = ap_fifo_oarg_74_din;
            assign tkeep[74] = {C_OUTPUT_FIFO_74_WIDTH/8{1'b1}};
            assign tstrb[74] = {C_OUTPUT_FIFO_74_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 75) begin
            assign dwconv_tready[75] = m_axis_fifo_75_tready;
            assign m_axis_fifo_75_tlast = dwconv_tlast[75];
            assign m_axis_fifo_75_tvalid = dwconv_tvalid[75];
            assign m_axis_fifo_75_tkeep = dwconv_tkeep[75][C_OUTPUT_FIFO_75_DMWIDTH/8-1:0];
            assign m_axis_fifo_75_tstrb = dwconv_tstrb[75][C_OUTPUT_FIFO_75_DMWIDTH/8-1:0];
            assign m_axis_fifo_75_tdata = dwconv_tdata[75][C_OUTPUT_FIFO_75_DMWIDTH-1:0];
            assign ap_fifo_oarg_75_full_n = full[75];
            assign write[75] = ap_fifo_oarg_75_write;
            assign din[75][C_OUTPUT_FIFO_75_WIDTH-1:0] = ap_fifo_oarg_75_din;
            assign tkeep[75] = {C_OUTPUT_FIFO_75_WIDTH/8{1'b1}};
            assign tstrb[75] = {C_OUTPUT_FIFO_75_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 76) begin
            assign dwconv_tready[76] = m_axis_fifo_76_tready;
            assign m_axis_fifo_76_tlast = dwconv_tlast[76];
            assign m_axis_fifo_76_tvalid = dwconv_tvalid[76];
            assign m_axis_fifo_76_tkeep = dwconv_tkeep[76][C_OUTPUT_FIFO_76_DMWIDTH/8-1:0];
            assign m_axis_fifo_76_tstrb = dwconv_tstrb[76][C_OUTPUT_FIFO_76_DMWIDTH/8-1:0];
            assign m_axis_fifo_76_tdata = dwconv_tdata[76][C_OUTPUT_FIFO_76_DMWIDTH-1:0];
            assign ap_fifo_oarg_76_full_n = full[76];
            assign write[76] = ap_fifo_oarg_76_write;
            assign din[76][C_OUTPUT_FIFO_76_WIDTH-1:0] = ap_fifo_oarg_76_din;
            assign tkeep[76] = {C_OUTPUT_FIFO_76_WIDTH/8{1'b1}};
            assign tstrb[76] = {C_OUTPUT_FIFO_76_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 77) begin
            assign dwconv_tready[77] = m_axis_fifo_77_tready;
            assign m_axis_fifo_77_tlast = dwconv_tlast[77];
            assign m_axis_fifo_77_tvalid = dwconv_tvalid[77];
            assign m_axis_fifo_77_tkeep = dwconv_tkeep[77][C_OUTPUT_FIFO_77_DMWIDTH/8-1:0];
            assign m_axis_fifo_77_tstrb = dwconv_tstrb[77][C_OUTPUT_FIFO_77_DMWIDTH/8-1:0];
            assign m_axis_fifo_77_tdata = dwconv_tdata[77][C_OUTPUT_FIFO_77_DMWIDTH-1:0];
            assign ap_fifo_oarg_77_full_n = full[77];
            assign write[77] = ap_fifo_oarg_77_write;
            assign din[77][C_OUTPUT_FIFO_77_WIDTH-1:0] = ap_fifo_oarg_77_din;
            assign tkeep[77] = {C_OUTPUT_FIFO_77_WIDTH/8{1'b1}};
            assign tstrb[77] = {C_OUTPUT_FIFO_77_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 78) begin
            assign dwconv_tready[78] = m_axis_fifo_78_tready;
            assign m_axis_fifo_78_tlast = dwconv_tlast[78];
            assign m_axis_fifo_78_tvalid = dwconv_tvalid[78];
            assign m_axis_fifo_78_tkeep = dwconv_tkeep[78][C_OUTPUT_FIFO_78_DMWIDTH/8-1:0];
            assign m_axis_fifo_78_tstrb = dwconv_tstrb[78][C_OUTPUT_FIFO_78_DMWIDTH/8-1:0];
            assign m_axis_fifo_78_tdata = dwconv_tdata[78][C_OUTPUT_FIFO_78_DMWIDTH-1:0];
            assign ap_fifo_oarg_78_full_n = full[78];
            assign write[78] = ap_fifo_oarg_78_write;
            assign din[78][C_OUTPUT_FIFO_78_WIDTH-1:0] = ap_fifo_oarg_78_din;
            assign tkeep[78] = {C_OUTPUT_FIFO_78_WIDTH/8{1'b1}};
            assign tstrb[78] = {C_OUTPUT_FIFO_78_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 79) begin
            assign dwconv_tready[79] = m_axis_fifo_79_tready;
            assign m_axis_fifo_79_tlast = dwconv_tlast[79];
            assign m_axis_fifo_79_tvalid = dwconv_tvalid[79];
            assign m_axis_fifo_79_tkeep = dwconv_tkeep[79][C_OUTPUT_FIFO_79_DMWIDTH/8-1:0];
            assign m_axis_fifo_79_tstrb = dwconv_tstrb[79][C_OUTPUT_FIFO_79_DMWIDTH/8-1:0];
            assign m_axis_fifo_79_tdata = dwconv_tdata[79][C_OUTPUT_FIFO_79_DMWIDTH-1:0];
            assign ap_fifo_oarg_79_full_n = full[79];
            assign write[79] = ap_fifo_oarg_79_write;
            assign din[79][C_OUTPUT_FIFO_79_WIDTH-1:0] = ap_fifo_oarg_79_din;
            assign tkeep[79] = {C_OUTPUT_FIFO_79_WIDTH/8{1'b1}};
            assign tstrb[79] = {C_OUTPUT_FIFO_79_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 80) begin
            assign dwconv_tready[80] = m_axis_fifo_80_tready;
            assign m_axis_fifo_80_tlast = dwconv_tlast[80];
            assign m_axis_fifo_80_tvalid = dwconv_tvalid[80];
            assign m_axis_fifo_80_tkeep = dwconv_tkeep[80][C_OUTPUT_FIFO_80_DMWIDTH/8-1:0];
            assign m_axis_fifo_80_tstrb = dwconv_tstrb[80][C_OUTPUT_FIFO_80_DMWIDTH/8-1:0];
            assign m_axis_fifo_80_tdata = dwconv_tdata[80][C_OUTPUT_FIFO_80_DMWIDTH-1:0];
            assign ap_fifo_oarg_80_full_n = full[80];
            assign write[80] = ap_fifo_oarg_80_write;
            assign din[80][C_OUTPUT_FIFO_80_WIDTH-1:0] = ap_fifo_oarg_80_din;
            assign tkeep[80] = {C_OUTPUT_FIFO_80_WIDTH/8{1'b1}};
            assign tstrb[80] = {C_OUTPUT_FIFO_80_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 81) begin
            assign dwconv_tready[81] = m_axis_fifo_81_tready;
            assign m_axis_fifo_81_tlast = dwconv_tlast[81];
            assign m_axis_fifo_81_tvalid = dwconv_tvalid[81];
            assign m_axis_fifo_81_tkeep = dwconv_tkeep[81][C_OUTPUT_FIFO_81_DMWIDTH/8-1:0];
            assign m_axis_fifo_81_tstrb = dwconv_tstrb[81][C_OUTPUT_FIFO_81_DMWIDTH/8-1:0];
            assign m_axis_fifo_81_tdata = dwconv_tdata[81][C_OUTPUT_FIFO_81_DMWIDTH-1:0];
            assign ap_fifo_oarg_81_full_n = full[81];
            assign write[81] = ap_fifo_oarg_81_write;
            assign din[81][C_OUTPUT_FIFO_81_WIDTH-1:0] = ap_fifo_oarg_81_din;
            assign tkeep[81] = {C_OUTPUT_FIFO_81_WIDTH/8{1'b1}};
            assign tstrb[81] = {C_OUTPUT_FIFO_81_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 82) begin
            assign dwconv_tready[82] = m_axis_fifo_82_tready;
            assign m_axis_fifo_82_tlast = dwconv_tlast[82];
            assign m_axis_fifo_82_tvalid = dwconv_tvalid[82];
            assign m_axis_fifo_82_tkeep = dwconv_tkeep[82][C_OUTPUT_FIFO_82_DMWIDTH/8-1:0];
            assign m_axis_fifo_82_tstrb = dwconv_tstrb[82][C_OUTPUT_FIFO_82_DMWIDTH/8-1:0];
            assign m_axis_fifo_82_tdata = dwconv_tdata[82][C_OUTPUT_FIFO_82_DMWIDTH-1:0];
            assign ap_fifo_oarg_82_full_n = full[82];
            assign write[82] = ap_fifo_oarg_82_write;
            assign din[82][C_OUTPUT_FIFO_82_WIDTH-1:0] = ap_fifo_oarg_82_din;
            assign tkeep[82] = {C_OUTPUT_FIFO_82_WIDTH/8{1'b1}};
            assign tstrb[82] = {C_OUTPUT_FIFO_82_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 83) begin
            assign dwconv_tready[83] = m_axis_fifo_83_tready;
            assign m_axis_fifo_83_tlast = dwconv_tlast[83];
            assign m_axis_fifo_83_tvalid = dwconv_tvalid[83];
            assign m_axis_fifo_83_tkeep = dwconv_tkeep[83][C_OUTPUT_FIFO_83_DMWIDTH/8-1:0];
            assign m_axis_fifo_83_tstrb = dwconv_tstrb[83][C_OUTPUT_FIFO_83_DMWIDTH/8-1:0];
            assign m_axis_fifo_83_tdata = dwconv_tdata[83][C_OUTPUT_FIFO_83_DMWIDTH-1:0];
            assign ap_fifo_oarg_83_full_n = full[83];
            assign write[83] = ap_fifo_oarg_83_write;
            assign din[83][C_OUTPUT_FIFO_83_WIDTH-1:0] = ap_fifo_oarg_83_din;
            assign tkeep[83] = {C_OUTPUT_FIFO_83_WIDTH/8{1'b1}};
            assign tstrb[83] = {C_OUTPUT_FIFO_83_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 84) begin
            assign dwconv_tready[84] = m_axis_fifo_84_tready;
            assign m_axis_fifo_84_tlast = dwconv_tlast[84];
            assign m_axis_fifo_84_tvalid = dwconv_tvalid[84];
            assign m_axis_fifo_84_tkeep = dwconv_tkeep[84][C_OUTPUT_FIFO_84_DMWIDTH/8-1:0];
            assign m_axis_fifo_84_tstrb = dwconv_tstrb[84][C_OUTPUT_FIFO_84_DMWIDTH/8-1:0];
            assign m_axis_fifo_84_tdata = dwconv_tdata[84][C_OUTPUT_FIFO_84_DMWIDTH-1:0];
            assign ap_fifo_oarg_84_full_n = full[84];
            assign write[84] = ap_fifo_oarg_84_write;
            assign din[84][C_OUTPUT_FIFO_84_WIDTH-1:0] = ap_fifo_oarg_84_din;
            assign tkeep[84] = {C_OUTPUT_FIFO_84_WIDTH/8{1'b1}};
            assign tstrb[84] = {C_OUTPUT_FIFO_84_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 85) begin
            assign dwconv_tready[85] = m_axis_fifo_85_tready;
            assign m_axis_fifo_85_tlast = dwconv_tlast[85];
            assign m_axis_fifo_85_tvalid = dwconv_tvalid[85];
            assign m_axis_fifo_85_tkeep = dwconv_tkeep[85][C_OUTPUT_FIFO_85_DMWIDTH/8-1:0];
            assign m_axis_fifo_85_tstrb = dwconv_tstrb[85][C_OUTPUT_FIFO_85_DMWIDTH/8-1:0];
            assign m_axis_fifo_85_tdata = dwconv_tdata[85][C_OUTPUT_FIFO_85_DMWIDTH-1:0];
            assign ap_fifo_oarg_85_full_n = full[85];
            assign write[85] = ap_fifo_oarg_85_write;
            assign din[85][C_OUTPUT_FIFO_85_WIDTH-1:0] = ap_fifo_oarg_85_din;
            assign tkeep[85] = {C_OUTPUT_FIFO_85_WIDTH/8{1'b1}};
            assign tstrb[85] = {C_OUTPUT_FIFO_85_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 86) begin
            assign dwconv_tready[86] = m_axis_fifo_86_tready;
            assign m_axis_fifo_86_tlast = dwconv_tlast[86];
            assign m_axis_fifo_86_tvalid = dwconv_tvalid[86];
            assign m_axis_fifo_86_tkeep = dwconv_tkeep[86][C_OUTPUT_FIFO_86_DMWIDTH/8-1:0];
            assign m_axis_fifo_86_tstrb = dwconv_tstrb[86][C_OUTPUT_FIFO_86_DMWIDTH/8-1:0];
            assign m_axis_fifo_86_tdata = dwconv_tdata[86][C_OUTPUT_FIFO_86_DMWIDTH-1:0];
            assign ap_fifo_oarg_86_full_n = full[86];
            assign write[86] = ap_fifo_oarg_86_write;
            assign din[86][C_OUTPUT_FIFO_86_WIDTH-1:0] = ap_fifo_oarg_86_din;
            assign tkeep[86] = {C_OUTPUT_FIFO_86_WIDTH/8{1'b1}};
            assign tstrb[86] = {C_OUTPUT_FIFO_86_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 87) begin
            assign dwconv_tready[87] = m_axis_fifo_87_tready;
            assign m_axis_fifo_87_tlast = dwconv_tlast[87];
            assign m_axis_fifo_87_tvalid = dwconv_tvalid[87];
            assign m_axis_fifo_87_tkeep = dwconv_tkeep[87][C_OUTPUT_FIFO_87_DMWIDTH/8-1:0];
            assign m_axis_fifo_87_tstrb = dwconv_tstrb[87][C_OUTPUT_FIFO_87_DMWIDTH/8-1:0];
            assign m_axis_fifo_87_tdata = dwconv_tdata[87][C_OUTPUT_FIFO_87_DMWIDTH-1:0];
            assign ap_fifo_oarg_87_full_n = full[87];
            assign write[87] = ap_fifo_oarg_87_write;
            assign din[87][C_OUTPUT_FIFO_87_WIDTH-1:0] = ap_fifo_oarg_87_din;
            assign tkeep[87] = {C_OUTPUT_FIFO_87_WIDTH/8{1'b1}};
            assign tstrb[87] = {C_OUTPUT_FIFO_87_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 88) begin
            assign dwconv_tready[88] = m_axis_fifo_88_tready;
            assign m_axis_fifo_88_tlast = dwconv_tlast[88];
            assign m_axis_fifo_88_tvalid = dwconv_tvalid[88];
            assign m_axis_fifo_88_tkeep = dwconv_tkeep[88][C_OUTPUT_FIFO_88_DMWIDTH/8-1:0];
            assign m_axis_fifo_88_tstrb = dwconv_tstrb[88][C_OUTPUT_FIFO_88_DMWIDTH/8-1:0];
            assign m_axis_fifo_88_tdata = dwconv_tdata[88][C_OUTPUT_FIFO_88_DMWIDTH-1:0];
            assign ap_fifo_oarg_88_full_n = full[88];
            assign write[88] = ap_fifo_oarg_88_write;
            assign din[88][C_OUTPUT_FIFO_88_WIDTH-1:0] = ap_fifo_oarg_88_din;
            assign tkeep[88] = {C_OUTPUT_FIFO_88_WIDTH/8{1'b1}};
            assign tstrb[88] = {C_OUTPUT_FIFO_88_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 89) begin
            assign dwconv_tready[89] = m_axis_fifo_89_tready;
            assign m_axis_fifo_89_tlast = dwconv_tlast[89];
            assign m_axis_fifo_89_tvalid = dwconv_tvalid[89];
            assign m_axis_fifo_89_tkeep = dwconv_tkeep[89][C_OUTPUT_FIFO_89_DMWIDTH/8-1:0];
            assign m_axis_fifo_89_tstrb = dwconv_tstrb[89][C_OUTPUT_FIFO_89_DMWIDTH/8-1:0];
            assign m_axis_fifo_89_tdata = dwconv_tdata[89][C_OUTPUT_FIFO_89_DMWIDTH-1:0];
            assign ap_fifo_oarg_89_full_n = full[89];
            assign write[89] = ap_fifo_oarg_89_write;
            assign din[89][C_OUTPUT_FIFO_89_WIDTH-1:0] = ap_fifo_oarg_89_din;
            assign tkeep[89] = {C_OUTPUT_FIFO_89_WIDTH/8{1'b1}};
            assign tstrb[89] = {C_OUTPUT_FIFO_89_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 90) begin
            assign dwconv_tready[90] = m_axis_fifo_90_tready;
            assign m_axis_fifo_90_tlast = dwconv_tlast[90];
            assign m_axis_fifo_90_tvalid = dwconv_tvalid[90];
            assign m_axis_fifo_90_tkeep = dwconv_tkeep[90][C_OUTPUT_FIFO_90_DMWIDTH/8-1:0];
            assign m_axis_fifo_90_tstrb = dwconv_tstrb[90][C_OUTPUT_FIFO_90_DMWIDTH/8-1:0];
            assign m_axis_fifo_90_tdata = dwconv_tdata[90][C_OUTPUT_FIFO_90_DMWIDTH-1:0];
            assign ap_fifo_oarg_90_full_n = full[90];
            assign write[90] = ap_fifo_oarg_90_write;
            assign din[90][C_OUTPUT_FIFO_90_WIDTH-1:0] = ap_fifo_oarg_90_din;
            assign tkeep[90] = {C_OUTPUT_FIFO_90_WIDTH/8{1'b1}};
            assign tstrb[90] = {C_OUTPUT_FIFO_90_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 91) begin
            assign dwconv_tready[91] = m_axis_fifo_91_tready;
            assign m_axis_fifo_91_tlast = dwconv_tlast[91];
            assign m_axis_fifo_91_tvalid = dwconv_tvalid[91];
            assign m_axis_fifo_91_tkeep = dwconv_tkeep[91][C_OUTPUT_FIFO_91_DMWIDTH/8-1:0];
            assign m_axis_fifo_91_tstrb = dwconv_tstrb[91][C_OUTPUT_FIFO_91_DMWIDTH/8-1:0];
            assign m_axis_fifo_91_tdata = dwconv_tdata[91][C_OUTPUT_FIFO_91_DMWIDTH-1:0];
            assign ap_fifo_oarg_91_full_n = full[91];
            assign write[91] = ap_fifo_oarg_91_write;
            assign din[91][C_OUTPUT_FIFO_91_WIDTH-1:0] = ap_fifo_oarg_91_din;
            assign tkeep[91] = {C_OUTPUT_FIFO_91_WIDTH/8{1'b1}};
            assign tstrb[91] = {C_OUTPUT_FIFO_91_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 92) begin
            assign dwconv_tready[92] = m_axis_fifo_92_tready;
            assign m_axis_fifo_92_tlast = dwconv_tlast[92];
            assign m_axis_fifo_92_tvalid = dwconv_tvalid[92];
            assign m_axis_fifo_92_tkeep = dwconv_tkeep[92][C_OUTPUT_FIFO_92_DMWIDTH/8-1:0];
            assign m_axis_fifo_92_tstrb = dwconv_tstrb[92][C_OUTPUT_FIFO_92_DMWIDTH/8-1:0];
            assign m_axis_fifo_92_tdata = dwconv_tdata[92][C_OUTPUT_FIFO_92_DMWIDTH-1:0];
            assign ap_fifo_oarg_92_full_n = full[92];
            assign write[92] = ap_fifo_oarg_92_write;
            assign din[92][C_OUTPUT_FIFO_92_WIDTH-1:0] = ap_fifo_oarg_92_din;
            assign tkeep[92] = {C_OUTPUT_FIFO_92_WIDTH/8{1'b1}};
            assign tstrb[92] = {C_OUTPUT_FIFO_92_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 93) begin
            assign dwconv_tready[93] = m_axis_fifo_93_tready;
            assign m_axis_fifo_93_tlast = dwconv_tlast[93];
            assign m_axis_fifo_93_tvalid = dwconv_tvalid[93];
            assign m_axis_fifo_93_tkeep = dwconv_tkeep[93][C_OUTPUT_FIFO_93_DMWIDTH/8-1:0];
            assign m_axis_fifo_93_tstrb = dwconv_tstrb[93][C_OUTPUT_FIFO_93_DMWIDTH/8-1:0];
            assign m_axis_fifo_93_tdata = dwconv_tdata[93][C_OUTPUT_FIFO_93_DMWIDTH-1:0];
            assign ap_fifo_oarg_93_full_n = full[93];
            assign write[93] = ap_fifo_oarg_93_write;
            assign din[93][C_OUTPUT_FIFO_93_WIDTH-1:0] = ap_fifo_oarg_93_din;
            assign tkeep[93] = {C_OUTPUT_FIFO_93_WIDTH/8{1'b1}};
            assign tstrb[93] = {C_OUTPUT_FIFO_93_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 94) begin
            assign dwconv_tready[94] = m_axis_fifo_94_tready;
            assign m_axis_fifo_94_tlast = dwconv_tlast[94];
            assign m_axis_fifo_94_tvalid = dwconv_tvalid[94];
            assign m_axis_fifo_94_tkeep = dwconv_tkeep[94][C_OUTPUT_FIFO_94_DMWIDTH/8-1:0];
            assign m_axis_fifo_94_tstrb = dwconv_tstrb[94][C_OUTPUT_FIFO_94_DMWIDTH/8-1:0];
            assign m_axis_fifo_94_tdata = dwconv_tdata[94][C_OUTPUT_FIFO_94_DMWIDTH-1:0];
            assign ap_fifo_oarg_94_full_n = full[94];
            assign write[94] = ap_fifo_oarg_94_write;
            assign din[94][C_OUTPUT_FIFO_94_WIDTH-1:0] = ap_fifo_oarg_94_din;
            assign tkeep[94] = {C_OUTPUT_FIFO_94_WIDTH/8{1'b1}};
            assign tstrb[94] = {C_OUTPUT_FIFO_94_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 95) begin
            assign dwconv_tready[95] = m_axis_fifo_95_tready;
            assign m_axis_fifo_95_tlast = dwconv_tlast[95];
            assign m_axis_fifo_95_tvalid = dwconv_tvalid[95];
            assign m_axis_fifo_95_tkeep = dwconv_tkeep[95][C_OUTPUT_FIFO_95_DMWIDTH/8-1:0];
            assign m_axis_fifo_95_tstrb = dwconv_tstrb[95][C_OUTPUT_FIFO_95_DMWIDTH/8-1:0];
            assign m_axis_fifo_95_tdata = dwconv_tdata[95][C_OUTPUT_FIFO_95_DMWIDTH-1:0];
            assign ap_fifo_oarg_95_full_n = full[95];
            assign write[95] = ap_fifo_oarg_95_write;
            assign din[95][C_OUTPUT_FIFO_95_WIDTH-1:0] = ap_fifo_oarg_95_din;
            assign tkeep[95] = {C_OUTPUT_FIFO_95_WIDTH/8{1'b1}};
            assign tstrb[95] = {C_OUTPUT_FIFO_95_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 96) begin
            assign dwconv_tready[96] = m_axis_fifo_96_tready;
            assign m_axis_fifo_96_tlast = dwconv_tlast[96];
            assign m_axis_fifo_96_tvalid = dwconv_tvalid[96];
            assign m_axis_fifo_96_tkeep = dwconv_tkeep[96][C_OUTPUT_FIFO_96_DMWIDTH/8-1:0];
            assign m_axis_fifo_96_tstrb = dwconv_tstrb[96][C_OUTPUT_FIFO_96_DMWIDTH/8-1:0];
            assign m_axis_fifo_96_tdata = dwconv_tdata[96][C_OUTPUT_FIFO_96_DMWIDTH-1:0];
            assign ap_fifo_oarg_96_full_n = full[96];
            assign write[96] = ap_fifo_oarg_96_write;
            assign din[96][C_OUTPUT_FIFO_96_WIDTH-1:0] = ap_fifo_oarg_96_din;
            assign tkeep[96] = {C_OUTPUT_FIFO_96_WIDTH/8{1'b1}};
            assign tstrb[96] = {C_OUTPUT_FIFO_96_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 97) begin
            assign dwconv_tready[97] = m_axis_fifo_97_tready;
            assign m_axis_fifo_97_tlast = dwconv_tlast[97];
            assign m_axis_fifo_97_tvalid = dwconv_tvalid[97];
            assign m_axis_fifo_97_tkeep = dwconv_tkeep[97][C_OUTPUT_FIFO_97_DMWIDTH/8-1:0];
            assign m_axis_fifo_97_tstrb = dwconv_tstrb[97][C_OUTPUT_FIFO_97_DMWIDTH/8-1:0];
            assign m_axis_fifo_97_tdata = dwconv_tdata[97][C_OUTPUT_FIFO_97_DMWIDTH-1:0];
            assign ap_fifo_oarg_97_full_n = full[97];
            assign write[97] = ap_fifo_oarg_97_write;
            assign din[97][C_OUTPUT_FIFO_97_WIDTH-1:0] = ap_fifo_oarg_97_din;
            assign tkeep[97] = {C_OUTPUT_FIFO_97_WIDTH/8{1'b1}};
            assign tstrb[97] = {C_OUTPUT_FIFO_97_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 98) begin
            assign dwconv_tready[98] = m_axis_fifo_98_tready;
            assign m_axis_fifo_98_tlast = dwconv_tlast[98];
            assign m_axis_fifo_98_tvalid = dwconv_tvalid[98];
            assign m_axis_fifo_98_tkeep = dwconv_tkeep[98][C_OUTPUT_FIFO_98_DMWIDTH/8-1:0];
            assign m_axis_fifo_98_tstrb = dwconv_tstrb[98][C_OUTPUT_FIFO_98_DMWIDTH/8-1:0];
            assign m_axis_fifo_98_tdata = dwconv_tdata[98][C_OUTPUT_FIFO_98_DMWIDTH-1:0];
            assign ap_fifo_oarg_98_full_n = full[98];
            assign write[98] = ap_fifo_oarg_98_write;
            assign din[98][C_OUTPUT_FIFO_98_WIDTH-1:0] = ap_fifo_oarg_98_din;
            assign tkeep[98] = {C_OUTPUT_FIFO_98_WIDTH/8{1'b1}};
            assign tstrb[98] = {C_OUTPUT_FIFO_98_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 99) begin
            assign dwconv_tready[99] = m_axis_fifo_99_tready;
            assign m_axis_fifo_99_tlast = dwconv_tlast[99];
            assign m_axis_fifo_99_tvalid = dwconv_tvalid[99];
            assign m_axis_fifo_99_tkeep = dwconv_tkeep[99][C_OUTPUT_FIFO_99_DMWIDTH/8-1:0];
            assign m_axis_fifo_99_tstrb = dwconv_tstrb[99][C_OUTPUT_FIFO_99_DMWIDTH/8-1:0];
            assign m_axis_fifo_99_tdata = dwconv_tdata[99][C_OUTPUT_FIFO_99_DMWIDTH-1:0];
            assign ap_fifo_oarg_99_full_n = full[99];
            assign write[99] = ap_fifo_oarg_99_write;
            assign din[99][C_OUTPUT_FIFO_99_WIDTH-1:0] = ap_fifo_oarg_99_din;
            assign tkeep[99] = {C_OUTPUT_FIFO_99_WIDTH/8{1'b1}};
            assign tstrb[99] = {C_OUTPUT_FIFO_99_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 100) begin
            assign dwconv_tready[100] = m_axis_fifo_100_tready;
            assign m_axis_fifo_100_tlast = dwconv_tlast[100];
            assign m_axis_fifo_100_tvalid = dwconv_tvalid[100];
            assign m_axis_fifo_100_tkeep = dwconv_tkeep[100][C_OUTPUT_FIFO_100_DMWIDTH/8-1:0];
            assign m_axis_fifo_100_tstrb = dwconv_tstrb[100][C_OUTPUT_FIFO_100_DMWIDTH/8-1:0];
            assign m_axis_fifo_100_tdata = dwconv_tdata[100][C_OUTPUT_FIFO_100_DMWIDTH-1:0];
            assign ap_fifo_oarg_100_full_n = full[100];
            assign write[100] = ap_fifo_oarg_100_write;
            assign din[100][C_OUTPUT_FIFO_100_WIDTH-1:0] = ap_fifo_oarg_100_din;
            assign tkeep[100] = {C_OUTPUT_FIFO_100_WIDTH/8{1'b1}};
            assign tstrb[100] = {C_OUTPUT_FIFO_100_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 101) begin
            assign dwconv_tready[101] = m_axis_fifo_101_tready;
            assign m_axis_fifo_101_tlast = dwconv_tlast[101];
            assign m_axis_fifo_101_tvalid = dwconv_tvalid[101];
            assign m_axis_fifo_101_tkeep = dwconv_tkeep[101][C_OUTPUT_FIFO_101_DMWIDTH/8-1:0];
            assign m_axis_fifo_101_tstrb = dwconv_tstrb[101][C_OUTPUT_FIFO_101_DMWIDTH/8-1:0];
            assign m_axis_fifo_101_tdata = dwconv_tdata[101][C_OUTPUT_FIFO_101_DMWIDTH-1:0];
            assign ap_fifo_oarg_101_full_n = full[101];
            assign write[101] = ap_fifo_oarg_101_write;
            assign din[101][C_OUTPUT_FIFO_101_WIDTH-1:0] = ap_fifo_oarg_101_din;
            assign tkeep[101] = {C_OUTPUT_FIFO_101_WIDTH/8{1'b1}};
            assign tstrb[101] = {C_OUTPUT_FIFO_101_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 102) begin
            assign dwconv_tready[102] = m_axis_fifo_102_tready;
            assign m_axis_fifo_102_tlast = dwconv_tlast[102];
            assign m_axis_fifo_102_tvalid = dwconv_tvalid[102];
            assign m_axis_fifo_102_tkeep = dwconv_tkeep[102][C_OUTPUT_FIFO_102_DMWIDTH/8-1:0];
            assign m_axis_fifo_102_tstrb = dwconv_tstrb[102][C_OUTPUT_FIFO_102_DMWIDTH/8-1:0];
            assign m_axis_fifo_102_tdata = dwconv_tdata[102][C_OUTPUT_FIFO_102_DMWIDTH-1:0];
            assign ap_fifo_oarg_102_full_n = full[102];
            assign write[102] = ap_fifo_oarg_102_write;
            assign din[102][C_OUTPUT_FIFO_102_WIDTH-1:0] = ap_fifo_oarg_102_din;
            assign tkeep[102] = {C_OUTPUT_FIFO_102_WIDTH/8{1'b1}};
            assign tstrb[102] = {C_OUTPUT_FIFO_102_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 103) begin
            assign dwconv_tready[103] = m_axis_fifo_103_tready;
            assign m_axis_fifo_103_tlast = dwconv_tlast[103];
            assign m_axis_fifo_103_tvalid = dwconv_tvalid[103];
            assign m_axis_fifo_103_tkeep = dwconv_tkeep[103][C_OUTPUT_FIFO_103_DMWIDTH/8-1:0];
            assign m_axis_fifo_103_tstrb = dwconv_tstrb[103][C_OUTPUT_FIFO_103_DMWIDTH/8-1:0];
            assign m_axis_fifo_103_tdata = dwconv_tdata[103][C_OUTPUT_FIFO_103_DMWIDTH-1:0];
            assign ap_fifo_oarg_103_full_n = full[103];
            assign write[103] = ap_fifo_oarg_103_write;
            assign din[103][C_OUTPUT_FIFO_103_WIDTH-1:0] = ap_fifo_oarg_103_din;
            assign tkeep[103] = {C_OUTPUT_FIFO_103_WIDTH/8{1'b1}};
            assign tstrb[103] = {C_OUTPUT_FIFO_103_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 104) begin
            assign dwconv_tready[104] = m_axis_fifo_104_tready;
            assign m_axis_fifo_104_tlast = dwconv_tlast[104];
            assign m_axis_fifo_104_tvalid = dwconv_tvalid[104];
            assign m_axis_fifo_104_tkeep = dwconv_tkeep[104][C_OUTPUT_FIFO_104_DMWIDTH/8-1:0];
            assign m_axis_fifo_104_tstrb = dwconv_tstrb[104][C_OUTPUT_FIFO_104_DMWIDTH/8-1:0];
            assign m_axis_fifo_104_tdata = dwconv_tdata[104][C_OUTPUT_FIFO_104_DMWIDTH-1:0];
            assign ap_fifo_oarg_104_full_n = full[104];
            assign write[104] = ap_fifo_oarg_104_write;
            assign din[104][C_OUTPUT_FIFO_104_WIDTH-1:0] = ap_fifo_oarg_104_din;
            assign tkeep[104] = {C_OUTPUT_FIFO_104_WIDTH/8{1'b1}};
            assign tstrb[104] = {C_OUTPUT_FIFO_104_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 105) begin
            assign dwconv_tready[105] = m_axis_fifo_105_tready;
            assign m_axis_fifo_105_tlast = dwconv_tlast[105];
            assign m_axis_fifo_105_tvalid = dwconv_tvalid[105];
            assign m_axis_fifo_105_tkeep = dwconv_tkeep[105][C_OUTPUT_FIFO_105_DMWIDTH/8-1:0];
            assign m_axis_fifo_105_tstrb = dwconv_tstrb[105][C_OUTPUT_FIFO_105_DMWIDTH/8-1:0];
            assign m_axis_fifo_105_tdata = dwconv_tdata[105][C_OUTPUT_FIFO_105_DMWIDTH-1:0];
            assign ap_fifo_oarg_105_full_n = full[105];
            assign write[105] = ap_fifo_oarg_105_write;
            assign din[105][C_OUTPUT_FIFO_105_WIDTH-1:0] = ap_fifo_oarg_105_din;
            assign tkeep[105] = {C_OUTPUT_FIFO_105_WIDTH/8{1'b1}};
            assign tstrb[105] = {C_OUTPUT_FIFO_105_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 106) begin
            assign dwconv_tready[106] = m_axis_fifo_106_tready;
            assign m_axis_fifo_106_tlast = dwconv_tlast[106];
            assign m_axis_fifo_106_tvalid = dwconv_tvalid[106];
            assign m_axis_fifo_106_tkeep = dwconv_tkeep[106][C_OUTPUT_FIFO_106_DMWIDTH/8-1:0];
            assign m_axis_fifo_106_tstrb = dwconv_tstrb[106][C_OUTPUT_FIFO_106_DMWIDTH/8-1:0];
            assign m_axis_fifo_106_tdata = dwconv_tdata[106][C_OUTPUT_FIFO_106_DMWIDTH-1:0];
            assign ap_fifo_oarg_106_full_n = full[106];
            assign write[106] = ap_fifo_oarg_106_write;
            assign din[106][C_OUTPUT_FIFO_106_WIDTH-1:0] = ap_fifo_oarg_106_din;
            assign tkeep[106] = {C_OUTPUT_FIFO_106_WIDTH/8{1'b1}};
            assign tstrb[106] = {C_OUTPUT_FIFO_106_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 107) begin
            assign dwconv_tready[107] = m_axis_fifo_107_tready;
            assign m_axis_fifo_107_tlast = dwconv_tlast[107];
            assign m_axis_fifo_107_tvalid = dwconv_tvalid[107];
            assign m_axis_fifo_107_tkeep = dwconv_tkeep[107][C_OUTPUT_FIFO_107_DMWIDTH/8-1:0];
            assign m_axis_fifo_107_tstrb = dwconv_tstrb[107][C_OUTPUT_FIFO_107_DMWIDTH/8-1:0];
            assign m_axis_fifo_107_tdata = dwconv_tdata[107][C_OUTPUT_FIFO_107_DMWIDTH-1:0];
            assign ap_fifo_oarg_107_full_n = full[107];
            assign write[107] = ap_fifo_oarg_107_write;
            assign din[107][C_OUTPUT_FIFO_107_WIDTH-1:0] = ap_fifo_oarg_107_din;
            assign tkeep[107] = {C_OUTPUT_FIFO_107_WIDTH/8{1'b1}};
            assign tstrb[107] = {C_OUTPUT_FIFO_107_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 108) begin
            assign dwconv_tready[108] = m_axis_fifo_108_tready;
            assign m_axis_fifo_108_tlast = dwconv_tlast[108];
            assign m_axis_fifo_108_tvalid = dwconv_tvalid[108];
            assign m_axis_fifo_108_tkeep = dwconv_tkeep[108][C_OUTPUT_FIFO_108_DMWIDTH/8-1:0];
            assign m_axis_fifo_108_tstrb = dwconv_tstrb[108][C_OUTPUT_FIFO_108_DMWIDTH/8-1:0];
            assign m_axis_fifo_108_tdata = dwconv_tdata[108][C_OUTPUT_FIFO_108_DMWIDTH-1:0];
            assign ap_fifo_oarg_108_full_n = full[108];
            assign write[108] = ap_fifo_oarg_108_write;
            assign din[108][C_OUTPUT_FIFO_108_WIDTH-1:0] = ap_fifo_oarg_108_din;
            assign tkeep[108] = {C_OUTPUT_FIFO_108_WIDTH/8{1'b1}};
            assign tstrb[108] = {C_OUTPUT_FIFO_108_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 109) begin
            assign dwconv_tready[109] = m_axis_fifo_109_tready;
            assign m_axis_fifo_109_tlast = dwconv_tlast[109];
            assign m_axis_fifo_109_tvalid = dwconv_tvalid[109];
            assign m_axis_fifo_109_tkeep = dwconv_tkeep[109][C_OUTPUT_FIFO_109_DMWIDTH/8-1:0];
            assign m_axis_fifo_109_tstrb = dwconv_tstrb[109][C_OUTPUT_FIFO_109_DMWIDTH/8-1:0];
            assign m_axis_fifo_109_tdata = dwconv_tdata[109][C_OUTPUT_FIFO_109_DMWIDTH-1:0];
            assign ap_fifo_oarg_109_full_n = full[109];
            assign write[109] = ap_fifo_oarg_109_write;
            assign din[109][C_OUTPUT_FIFO_109_WIDTH-1:0] = ap_fifo_oarg_109_din;
            assign tkeep[109] = {C_OUTPUT_FIFO_109_WIDTH/8{1'b1}};
            assign tstrb[109] = {C_OUTPUT_FIFO_109_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 110) begin
            assign dwconv_tready[110] = m_axis_fifo_110_tready;
            assign m_axis_fifo_110_tlast = dwconv_tlast[110];
            assign m_axis_fifo_110_tvalid = dwconv_tvalid[110];
            assign m_axis_fifo_110_tkeep = dwconv_tkeep[110][C_OUTPUT_FIFO_110_DMWIDTH/8-1:0];
            assign m_axis_fifo_110_tstrb = dwconv_tstrb[110][C_OUTPUT_FIFO_110_DMWIDTH/8-1:0];
            assign m_axis_fifo_110_tdata = dwconv_tdata[110][C_OUTPUT_FIFO_110_DMWIDTH-1:0];
            assign ap_fifo_oarg_110_full_n = full[110];
            assign write[110] = ap_fifo_oarg_110_write;
            assign din[110][C_OUTPUT_FIFO_110_WIDTH-1:0] = ap_fifo_oarg_110_din;
            assign tkeep[110] = {C_OUTPUT_FIFO_110_WIDTH/8{1'b1}};
            assign tstrb[110] = {C_OUTPUT_FIFO_110_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 111) begin
            assign dwconv_tready[111] = m_axis_fifo_111_tready;
            assign m_axis_fifo_111_tlast = dwconv_tlast[111];
            assign m_axis_fifo_111_tvalid = dwconv_tvalid[111];
            assign m_axis_fifo_111_tkeep = dwconv_tkeep[111][C_OUTPUT_FIFO_111_DMWIDTH/8-1:0];
            assign m_axis_fifo_111_tstrb = dwconv_tstrb[111][C_OUTPUT_FIFO_111_DMWIDTH/8-1:0];
            assign m_axis_fifo_111_tdata = dwconv_tdata[111][C_OUTPUT_FIFO_111_DMWIDTH-1:0];
            assign ap_fifo_oarg_111_full_n = full[111];
            assign write[111] = ap_fifo_oarg_111_write;
            assign din[111][C_OUTPUT_FIFO_111_WIDTH-1:0] = ap_fifo_oarg_111_din;
            assign tkeep[111] = {C_OUTPUT_FIFO_111_WIDTH/8{1'b1}};
            assign tstrb[111] = {C_OUTPUT_FIFO_111_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 112) begin
            assign dwconv_tready[112] = m_axis_fifo_112_tready;
            assign m_axis_fifo_112_tlast = dwconv_tlast[112];
            assign m_axis_fifo_112_tvalid = dwconv_tvalid[112];
            assign m_axis_fifo_112_tkeep = dwconv_tkeep[112][C_OUTPUT_FIFO_112_DMWIDTH/8-1:0];
            assign m_axis_fifo_112_tstrb = dwconv_tstrb[112][C_OUTPUT_FIFO_112_DMWIDTH/8-1:0];
            assign m_axis_fifo_112_tdata = dwconv_tdata[112][C_OUTPUT_FIFO_112_DMWIDTH-1:0];
            assign ap_fifo_oarg_112_full_n = full[112];
            assign write[112] = ap_fifo_oarg_112_write;
            assign din[112][C_OUTPUT_FIFO_112_WIDTH-1:0] = ap_fifo_oarg_112_din;
            assign tkeep[112] = {C_OUTPUT_FIFO_112_WIDTH/8{1'b1}};
            assign tstrb[112] = {C_OUTPUT_FIFO_112_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 113) begin
            assign dwconv_tready[113] = m_axis_fifo_113_tready;
            assign m_axis_fifo_113_tlast = dwconv_tlast[113];
            assign m_axis_fifo_113_tvalid = dwconv_tvalid[113];
            assign m_axis_fifo_113_tkeep = dwconv_tkeep[113][C_OUTPUT_FIFO_113_DMWIDTH/8-1:0];
            assign m_axis_fifo_113_tstrb = dwconv_tstrb[113][C_OUTPUT_FIFO_113_DMWIDTH/8-1:0];
            assign m_axis_fifo_113_tdata = dwconv_tdata[113][C_OUTPUT_FIFO_113_DMWIDTH-1:0];
            assign ap_fifo_oarg_113_full_n = full[113];
            assign write[113] = ap_fifo_oarg_113_write;
            assign din[113][C_OUTPUT_FIFO_113_WIDTH-1:0] = ap_fifo_oarg_113_din;
            assign tkeep[113] = {C_OUTPUT_FIFO_113_WIDTH/8{1'b1}};
            assign tstrb[113] = {C_OUTPUT_FIFO_113_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 114) begin
            assign dwconv_tready[114] = m_axis_fifo_114_tready;
            assign m_axis_fifo_114_tlast = dwconv_tlast[114];
            assign m_axis_fifo_114_tvalid = dwconv_tvalid[114];
            assign m_axis_fifo_114_tkeep = dwconv_tkeep[114][C_OUTPUT_FIFO_114_DMWIDTH/8-1:0];
            assign m_axis_fifo_114_tstrb = dwconv_tstrb[114][C_OUTPUT_FIFO_114_DMWIDTH/8-1:0];
            assign m_axis_fifo_114_tdata = dwconv_tdata[114][C_OUTPUT_FIFO_114_DMWIDTH-1:0];
            assign ap_fifo_oarg_114_full_n = full[114];
            assign write[114] = ap_fifo_oarg_114_write;
            assign din[114][C_OUTPUT_FIFO_114_WIDTH-1:0] = ap_fifo_oarg_114_din;
            assign tkeep[114] = {C_OUTPUT_FIFO_114_WIDTH/8{1'b1}};
            assign tstrb[114] = {C_OUTPUT_FIFO_114_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 115) begin
            assign dwconv_tready[115] = m_axis_fifo_115_tready;
            assign m_axis_fifo_115_tlast = dwconv_tlast[115];
            assign m_axis_fifo_115_tvalid = dwconv_tvalid[115];
            assign m_axis_fifo_115_tkeep = dwconv_tkeep[115][C_OUTPUT_FIFO_115_DMWIDTH/8-1:0];
            assign m_axis_fifo_115_tstrb = dwconv_tstrb[115][C_OUTPUT_FIFO_115_DMWIDTH/8-1:0];
            assign m_axis_fifo_115_tdata = dwconv_tdata[115][C_OUTPUT_FIFO_115_DMWIDTH-1:0];
            assign ap_fifo_oarg_115_full_n = full[115];
            assign write[115] = ap_fifo_oarg_115_write;
            assign din[115][C_OUTPUT_FIFO_115_WIDTH-1:0] = ap_fifo_oarg_115_din;
            assign tkeep[115] = {C_OUTPUT_FIFO_115_WIDTH/8{1'b1}};
            assign tstrb[115] = {C_OUTPUT_FIFO_115_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 116) begin
            assign dwconv_tready[116] = m_axis_fifo_116_tready;
            assign m_axis_fifo_116_tlast = dwconv_tlast[116];
            assign m_axis_fifo_116_tvalid = dwconv_tvalid[116];
            assign m_axis_fifo_116_tkeep = dwconv_tkeep[116][C_OUTPUT_FIFO_116_DMWIDTH/8-1:0];
            assign m_axis_fifo_116_tstrb = dwconv_tstrb[116][C_OUTPUT_FIFO_116_DMWIDTH/8-1:0];
            assign m_axis_fifo_116_tdata = dwconv_tdata[116][C_OUTPUT_FIFO_116_DMWIDTH-1:0];
            assign ap_fifo_oarg_116_full_n = full[116];
            assign write[116] = ap_fifo_oarg_116_write;
            assign din[116][C_OUTPUT_FIFO_116_WIDTH-1:0] = ap_fifo_oarg_116_din;
            assign tkeep[116] = {C_OUTPUT_FIFO_116_WIDTH/8{1'b1}};
            assign tstrb[116] = {C_OUTPUT_FIFO_116_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 117) begin
            assign dwconv_tready[117] = m_axis_fifo_117_tready;
            assign m_axis_fifo_117_tlast = dwconv_tlast[117];
            assign m_axis_fifo_117_tvalid = dwconv_tvalid[117];
            assign m_axis_fifo_117_tkeep = dwconv_tkeep[117][C_OUTPUT_FIFO_117_DMWIDTH/8-1:0];
            assign m_axis_fifo_117_tstrb = dwconv_tstrb[117][C_OUTPUT_FIFO_117_DMWIDTH/8-1:0];
            assign m_axis_fifo_117_tdata = dwconv_tdata[117][C_OUTPUT_FIFO_117_DMWIDTH-1:0];
            assign ap_fifo_oarg_117_full_n = full[117];
            assign write[117] = ap_fifo_oarg_117_write;
            assign din[117][C_OUTPUT_FIFO_117_WIDTH-1:0] = ap_fifo_oarg_117_din;
            assign tkeep[117] = {C_OUTPUT_FIFO_117_WIDTH/8{1'b1}};
            assign tstrb[117] = {C_OUTPUT_FIFO_117_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 118) begin
            assign dwconv_tready[118] = m_axis_fifo_118_tready;
            assign m_axis_fifo_118_tlast = dwconv_tlast[118];
            assign m_axis_fifo_118_tvalid = dwconv_tvalid[118];
            assign m_axis_fifo_118_tkeep = dwconv_tkeep[118][C_OUTPUT_FIFO_118_DMWIDTH/8-1:0];
            assign m_axis_fifo_118_tstrb = dwconv_tstrb[118][C_OUTPUT_FIFO_118_DMWIDTH/8-1:0];
            assign m_axis_fifo_118_tdata = dwconv_tdata[118][C_OUTPUT_FIFO_118_DMWIDTH-1:0];
            assign ap_fifo_oarg_118_full_n = full[118];
            assign write[118] = ap_fifo_oarg_118_write;
            assign din[118][C_OUTPUT_FIFO_118_WIDTH-1:0] = ap_fifo_oarg_118_din;
            assign tkeep[118] = {C_OUTPUT_FIFO_118_WIDTH/8{1'b1}};
            assign tstrb[118] = {C_OUTPUT_FIFO_118_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 119) begin
            assign dwconv_tready[119] = m_axis_fifo_119_tready;
            assign m_axis_fifo_119_tlast = dwconv_tlast[119];
            assign m_axis_fifo_119_tvalid = dwconv_tvalid[119];
            assign m_axis_fifo_119_tkeep = dwconv_tkeep[119][C_OUTPUT_FIFO_119_DMWIDTH/8-1:0];
            assign m_axis_fifo_119_tstrb = dwconv_tstrb[119][C_OUTPUT_FIFO_119_DMWIDTH/8-1:0];
            assign m_axis_fifo_119_tdata = dwconv_tdata[119][C_OUTPUT_FIFO_119_DMWIDTH-1:0];
            assign ap_fifo_oarg_119_full_n = full[119];
            assign write[119] = ap_fifo_oarg_119_write;
            assign din[119][C_OUTPUT_FIFO_119_WIDTH-1:0] = ap_fifo_oarg_119_din;
            assign tkeep[119] = {C_OUTPUT_FIFO_119_WIDTH/8{1'b1}};
            assign tstrb[119] = {C_OUTPUT_FIFO_119_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 120) begin
            assign dwconv_tready[120] = m_axis_fifo_120_tready;
            assign m_axis_fifo_120_tlast = dwconv_tlast[120];
            assign m_axis_fifo_120_tvalid = dwconv_tvalid[120];
            assign m_axis_fifo_120_tkeep = dwconv_tkeep[120][C_OUTPUT_FIFO_120_DMWIDTH/8-1:0];
            assign m_axis_fifo_120_tstrb = dwconv_tstrb[120][C_OUTPUT_FIFO_120_DMWIDTH/8-1:0];
            assign m_axis_fifo_120_tdata = dwconv_tdata[120][C_OUTPUT_FIFO_120_DMWIDTH-1:0];
            assign ap_fifo_oarg_120_full_n = full[120];
            assign write[120] = ap_fifo_oarg_120_write;
            assign din[120][C_OUTPUT_FIFO_120_WIDTH-1:0] = ap_fifo_oarg_120_din;
            assign tkeep[120] = {C_OUTPUT_FIFO_120_WIDTH/8{1'b1}};
            assign tstrb[120] = {C_OUTPUT_FIFO_120_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 121) begin
            assign dwconv_tready[121] = m_axis_fifo_121_tready;
            assign m_axis_fifo_121_tlast = dwconv_tlast[121];
            assign m_axis_fifo_121_tvalid = dwconv_tvalid[121];
            assign m_axis_fifo_121_tkeep = dwconv_tkeep[121][C_OUTPUT_FIFO_121_DMWIDTH/8-1:0];
            assign m_axis_fifo_121_tstrb = dwconv_tstrb[121][C_OUTPUT_FIFO_121_DMWIDTH/8-1:0];
            assign m_axis_fifo_121_tdata = dwconv_tdata[121][C_OUTPUT_FIFO_121_DMWIDTH-1:0];
            assign ap_fifo_oarg_121_full_n = full[121];
            assign write[121] = ap_fifo_oarg_121_write;
            assign din[121][C_OUTPUT_FIFO_121_WIDTH-1:0] = ap_fifo_oarg_121_din;
            assign tkeep[121] = {C_OUTPUT_FIFO_121_WIDTH/8{1'b1}};
            assign tstrb[121] = {C_OUTPUT_FIFO_121_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 122) begin
            assign dwconv_tready[122] = m_axis_fifo_122_tready;
            assign m_axis_fifo_122_tlast = dwconv_tlast[122];
            assign m_axis_fifo_122_tvalid = dwconv_tvalid[122];
            assign m_axis_fifo_122_tkeep = dwconv_tkeep[122][C_OUTPUT_FIFO_122_DMWIDTH/8-1:0];
            assign m_axis_fifo_122_tstrb = dwconv_tstrb[122][C_OUTPUT_FIFO_122_DMWIDTH/8-1:0];
            assign m_axis_fifo_122_tdata = dwconv_tdata[122][C_OUTPUT_FIFO_122_DMWIDTH-1:0];
            assign ap_fifo_oarg_122_full_n = full[122];
            assign write[122] = ap_fifo_oarg_122_write;
            assign din[122][C_OUTPUT_FIFO_122_WIDTH-1:0] = ap_fifo_oarg_122_din;
            assign tkeep[122] = {C_OUTPUT_FIFO_122_WIDTH/8{1'b1}};
            assign tstrb[122] = {C_OUTPUT_FIFO_122_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 123) begin
            assign dwconv_tready[123] = m_axis_fifo_123_tready;
            assign m_axis_fifo_123_tlast = dwconv_tlast[123];
            assign m_axis_fifo_123_tvalid = dwconv_tvalid[123];
            assign m_axis_fifo_123_tkeep = dwconv_tkeep[123][C_OUTPUT_FIFO_123_DMWIDTH/8-1:0];
            assign m_axis_fifo_123_tstrb = dwconv_tstrb[123][C_OUTPUT_FIFO_123_DMWIDTH/8-1:0];
            assign m_axis_fifo_123_tdata = dwconv_tdata[123][C_OUTPUT_FIFO_123_DMWIDTH-1:0];
            assign ap_fifo_oarg_123_full_n = full[123];
            assign write[123] = ap_fifo_oarg_123_write;
            assign din[123][C_OUTPUT_FIFO_123_WIDTH-1:0] = ap_fifo_oarg_123_din;
            assign tkeep[123] = {C_OUTPUT_FIFO_123_WIDTH/8{1'b1}};
            assign tstrb[123] = {C_OUTPUT_FIFO_123_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 124) begin
            assign dwconv_tready[124] = m_axis_fifo_124_tready;
            assign m_axis_fifo_124_tlast = dwconv_tlast[124];
            assign m_axis_fifo_124_tvalid = dwconv_tvalid[124];
            assign m_axis_fifo_124_tkeep = dwconv_tkeep[124][C_OUTPUT_FIFO_124_DMWIDTH/8-1:0];
            assign m_axis_fifo_124_tstrb = dwconv_tstrb[124][C_OUTPUT_FIFO_124_DMWIDTH/8-1:0];
            assign m_axis_fifo_124_tdata = dwconv_tdata[124][C_OUTPUT_FIFO_124_DMWIDTH-1:0];
            assign ap_fifo_oarg_124_full_n = full[124];
            assign write[124] = ap_fifo_oarg_124_write;
            assign din[124][C_OUTPUT_FIFO_124_WIDTH-1:0] = ap_fifo_oarg_124_din;
            assign tkeep[124] = {C_OUTPUT_FIFO_124_WIDTH/8{1'b1}};
            assign tstrb[124] = {C_OUTPUT_FIFO_124_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 125) begin
            assign dwconv_tready[125] = m_axis_fifo_125_tready;
            assign m_axis_fifo_125_tlast = dwconv_tlast[125];
            assign m_axis_fifo_125_tvalid = dwconv_tvalid[125];
            assign m_axis_fifo_125_tkeep = dwconv_tkeep[125][C_OUTPUT_FIFO_125_DMWIDTH/8-1:0];
            assign m_axis_fifo_125_tstrb = dwconv_tstrb[125][C_OUTPUT_FIFO_125_DMWIDTH/8-1:0];
            assign m_axis_fifo_125_tdata = dwconv_tdata[125][C_OUTPUT_FIFO_125_DMWIDTH-1:0];
            assign ap_fifo_oarg_125_full_n = full[125];
            assign write[125] = ap_fifo_oarg_125_write;
            assign din[125][C_OUTPUT_FIFO_125_WIDTH-1:0] = ap_fifo_oarg_125_din;
            assign tkeep[125] = {C_OUTPUT_FIFO_125_WIDTH/8{1'b1}};
            assign tstrb[125] = {C_OUTPUT_FIFO_125_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 126) begin
            assign dwconv_tready[126] = m_axis_fifo_126_tready;
            assign m_axis_fifo_126_tlast = dwconv_tlast[126];
            assign m_axis_fifo_126_tvalid = dwconv_tvalid[126];
            assign m_axis_fifo_126_tkeep = dwconv_tkeep[126][C_OUTPUT_FIFO_126_DMWIDTH/8-1:0];
            assign m_axis_fifo_126_tstrb = dwconv_tstrb[126][C_OUTPUT_FIFO_126_DMWIDTH/8-1:0];
            assign m_axis_fifo_126_tdata = dwconv_tdata[126][C_OUTPUT_FIFO_126_DMWIDTH-1:0];
            assign ap_fifo_oarg_126_full_n = full[126];
            assign write[126] = ap_fifo_oarg_126_write;
            assign din[126][C_OUTPUT_FIFO_126_WIDTH-1:0] = ap_fifo_oarg_126_din;
            assign tkeep[126] = {C_OUTPUT_FIFO_126_WIDTH/8{1'b1}};
            assign tstrb[126] = {C_OUTPUT_FIFO_126_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_FIFOs > 127) begin
            assign dwconv_tready[127] = m_axis_fifo_127_tready;
            assign m_axis_fifo_127_tlast = dwconv_tlast[127];
            assign m_axis_fifo_127_tvalid = dwconv_tvalid[127];
            assign m_axis_fifo_127_tkeep = dwconv_tkeep[127][C_OUTPUT_FIFO_127_DMWIDTH/8-1:0];
            assign m_axis_fifo_127_tstrb = dwconv_tstrb[127][C_OUTPUT_FIFO_127_DMWIDTH/8-1:0];
            assign m_axis_fifo_127_tdata = dwconv_tdata[127][C_OUTPUT_FIFO_127_DMWIDTH-1:0];
            assign ap_fifo_oarg_127_full_n = full[127];
            assign write[127] = ap_fifo_oarg_127_write;
            assign din[127][C_OUTPUT_FIFO_127_WIDTH-1:0] = ap_fifo_oarg_127_din;
            assign tkeep[127] = {C_OUTPUT_FIFO_127_WIDTH/8{1'b1}};
            assign tstrb[127] = {C_OUTPUT_FIFO_127_WIDTH/8{1'b1}};
        end
    endgenerate    
    
    //instantiate the axis2fifo modules
    genvar idx;
    generate
        for(idx=0; idx<C_NUM_OUTPUT_FIFOs; idx=idx+1) begin: OUT_FIFO_GEN
            fifo2axis #( 
                .DATA_WIDTH(C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx])
            ) fifo2axis_i (
                .ACC_CLK(acc_clk),
                .ARESETN(aresetn),
                .CTRL_ALLOW(out_fifo_allow),
                .CTRL_READY(out_fifo_ready[idx]),
                .CTRL_FINISHED(out_fifo_finished[idx]),
                .AXIS_TLAST(tlast[idx]),
                .AXIS_TVALID(tvalid[idx]),
                .AXIS_TDATA(tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .AXIS_TREADY(tready[idx]),
                .FIFO_FULL(full[idx]),
                .FIFO_DIN(din[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .FIFO_WRITE(write[idx])
            );
            
            //always use fifo
            axis_fifo #(
                .C_DATA_WIDTH(C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                .C_DATA_DEPTH(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx])
            ) axis_fifo_i (
                .aresetn(aresetn),
                .inclk(acc_clk),
                .in_tdata(tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .in_tlast(tlast[idx]),  
                .in_tvalid(tvalid[idx]),
                .in_tready(tready[idx]),
                .outclk(dm_clk), 
                .out_tdata(buf_tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .out_tready(buf_tready[idx]),
                .out_tvalid(buf_tvalid[idx]),
                .out_tlast(buf_tlast[idx])
            );
            
            //check if data width converter is needed
            if(C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx] != C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]) begin
                 axis_dwidth_converter_v1_1_9_axis_dwidth_converter #(
                    .C_S_AXIS_TDATA_WIDTH(C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_M_AXIS_TDATA_WIDTH(C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_AXIS_TID_WIDTH(1),
                    .C_AXIS_TDEST_WIDTH(1),
                    .C_S_AXIS_TUSER_WIDTH(1),
                    .C_M_AXIS_TUSER_WIDTH(1),
                    .C_AXIS_SIGNAL_SET(32'h1F)  //Enabled: TLAST, TKEEP, TSTRB, TDATA, TREADY
                ) data_width_conv_i (
                    .aclk(dm_clk),
                    .aresetn(aresetn),
                    .aclken(1),
                    .s_axis_tvalid(buf_tvalid[idx]),
                    .s_axis_tready(buf_tready[idx]),
                    .s_axis_tdata(buf_tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .s_axis_tstrb(tstrb[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tkeep(tkeep[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tlast(buf_tlast[idx]),
//                    .s_axis_tid(),
//                    .s_axis_tdest(),
//                    .s_axis_tuser(),
                    .m_axis_tvalid(dwconv_tvalid[idx]),
                    .m_axis_tready(dwconv_tready[idx]),
                    .m_axis_tdata(dwconv_tdata[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .m_axis_tstrb(dwconv_tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .m_axis_tkeep(dwconv_tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .m_axis_tlast(dwconv_tlast[idx])
//                    .m_axis_tid(),
//                    .m_axis_tdest(),
//                    .m_axis_tuser()
                );
            end
            else begin
                //if no data width converter, wire the input signals straight through
                assign dwconv_tlast[idx] = buf_tlast[idx];
                assign dwconv_tvalid[idx] = buf_tvalid[idx];
                assign buf_tready[idx] = dwconv_tready[idx];   //output
                assign dwconv_tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = buf_tdata[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
                assign dwconv_tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0] = tstrb[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0];
                assign dwconv_tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0] = tkeep[idx][C_OUTFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0];
            end
        end
    endgenerate
endmodule
