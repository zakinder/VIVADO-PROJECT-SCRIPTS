`timescale 1ns / 1ps

module top (
    //axi lite interface
    input s_axi_aclk,
    input s_axi_aresetn,
    input [31 : 0] S_AXI_AWADDR,
    input [2 : 0] S_AXI_AWPROT,
    input S_AXI_AWVALID,
    output S_AXI_AWREADY,
    input [31 : 0] S_AXI_WDATA,
    input [3 : 0] S_AXI_WSTRB,
    input S_AXI_WVALID,
    output S_AXI_WREADY,
    output [1 : 0] S_AXI_BRESP,
    output S_AXI_BVALID,
    input S_AXI_BREADY,
    input [31 : 0] S_AXI_ARADDR,
    input [2 : 0] S_AXI_ARPROT,
    input S_AXI_ARVALID,
    output S_AXI_ARREADY,
    output [31 : 0] S_AXI_RDATA,
    output [1 : 0] S_AXI_RRESP,
    output S_AXI_RVALID,
    input S_AXI_RREADY,
    //acc clock
    input aclk,
    input resetn,
    //acc interface
    output aresetn,
    output ap_start,
    input ap_idle,
    input ap_done,
    input ap_ready,
    output ap_continue,
    output ap_clk,
    //-----------------------------------------------------
    //input scalar ports
    output [C_INPUT_SCALAR_0_WIDTH-1:0] ap_iscalar_0_dout,
    output [C_INPUT_SCALAR_1_WIDTH-1:0] ap_iscalar_1_dout,
    output [C_INPUT_SCALAR_2_WIDTH-1:0] ap_iscalar_2_dout,
    output [C_INPUT_SCALAR_3_WIDTH-1:0] ap_iscalar_3_dout,
    output [C_INPUT_SCALAR_4_WIDTH-1:0] ap_iscalar_4_dout,
    output [C_INPUT_SCALAR_5_WIDTH-1:0] ap_iscalar_5_dout,
    output [C_INPUT_SCALAR_6_WIDTH-1:0] ap_iscalar_6_dout,
    output [C_INPUT_SCALAR_7_WIDTH-1:0] ap_iscalar_7_dout,
    output [C_INPUT_SCALAR_8_WIDTH-1:0] ap_iscalar_8_dout,
    output [C_INPUT_SCALAR_9_WIDTH-1:0] ap_iscalar_9_dout,
    output [C_INPUT_SCALAR_10_WIDTH-1:0] ap_iscalar_10_dout,
    output [C_INPUT_SCALAR_11_WIDTH-1:0] ap_iscalar_11_dout,
    output [C_INPUT_SCALAR_12_WIDTH-1:0] ap_iscalar_12_dout,
    output [C_INPUT_SCALAR_13_WIDTH-1:0] ap_iscalar_13_dout,
    output [C_INPUT_SCALAR_14_WIDTH-1:0] ap_iscalar_14_dout,
    output [C_INPUT_SCALAR_15_WIDTH-1:0] ap_iscalar_15_dout,
    output [C_INPUT_SCALAR_16_WIDTH-1:0] ap_iscalar_16_dout,
    output [C_INPUT_SCALAR_17_WIDTH-1:0] ap_iscalar_17_dout,
    output [C_INPUT_SCALAR_18_WIDTH-1:0] ap_iscalar_18_dout,
    output [C_INPUT_SCALAR_19_WIDTH-1:0] ap_iscalar_19_dout,
    output [C_INPUT_SCALAR_20_WIDTH-1:0] ap_iscalar_20_dout,
    output [C_INPUT_SCALAR_21_WIDTH-1:0] ap_iscalar_21_dout,
    output [C_INPUT_SCALAR_22_WIDTH-1:0] ap_iscalar_22_dout,
    output [C_INPUT_SCALAR_23_WIDTH-1:0] ap_iscalar_23_dout,
    output [C_INPUT_SCALAR_24_WIDTH-1:0] ap_iscalar_24_dout,
    output [C_INPUT_SCALAR_25_WIDTH-1:0] ap_iscalar_25_dout,
    output [C_INPUT_SCALAR_26_WIDTH-1:0] ap_iscalar_26_dout,
    output [C_INPUT_SCALAR_27_WIDTH-1:0] ap_iscalar_27_dout,
    output [C_INPUT_SCALAR_28_WIDTH-1:0] ap_iscalar_28_dout,
    output [C_INPUT_SCALAR_29_WIDTH-1:0] ap_iscalar_29_dout,
    output [C_INPUT_SCALAR_30_WIDTH-1:0] ap_iscalar_30_dout,
    output [C_INPUT_SCALAR_31_WIDTH-1:0] ap_iscalar_31_dout,
    output [C_INPUT_SCALAR_32_WIDTH-1:0] ap_iscalar_32_dout,
    output [C_INPUT_SCALAR_33_WIDTH-1:0] ap_iscalar_33_dout,
    output [C_INPUT_SCALAR_34_WIDTH-1:0] ap_iscalar_34_dout,
    output [C_INPUT_SCALAR_35_WIDTH-1:0] ap_iscalar_35_dout,
    output [C_INPUT_SCALAR_36_WIDTH-1:0] ap_iscalar_36_dout,
    output [C_INPUT_SCALAR_37_WIDTH-1:0] ap_iscalar_37_dout,
    output [C_INPUT_SCALAR_38_WIDTH-1:0] ap_iscalar_38_dout,
    output [C_INPUT_SCALAR_39_WIDTH-1:0] ap_iscalar_39_dout,
    output [C_INPUT_SCALAR_40_WIDTH-1:0] ap_iscalar_40_dout,
    output [C_INPUT_SCALAR_41_WIDTH-1:0] ap_iscalar_41_dout,
    output [C_INPUT_SCALAR_42_WIDTH-1:0] ap_iscalar_42_dout,
    output [C_INPUT_SCALAR_43_WIDTH-1:0] ap_iscalar_43_dout,
    output [C_INPUT_SCALAR_44_WIDTH-1:0] ap_iscalar_44_dout,
    output [C_INPUT_SCALAR_45_WIDTH-1:0] ap_iscalar_45_dout,
    output [C_INPUT_SCALAR_46_WIDTH-1:0] ap_iscalar_46_dout,
    output [C_INPUT_SCALAR_47_WIDTH-1:0] ap_iscalar_47_dout,
    output [C_INPUT_SCALAR_48_WIDTH-1:0] ap_iscalar_48_dout,
    output [C_INPUT_SCALAR_49_WIDTH-1:0] ap_iscalar_49_dout,
    output [C_INPUT_SCALAR_50_WIDTH-1:0] ap_iscalar_50_dout,
    output [C_INPUT_SCALAR_51_WIDTH-1:0] ap_iscalar_51_dout,
    output [C_INPUT_SCALAR_52_WIDTH-1:0] ap_iscalar_52_dout,
    output [C_INPUT_SCALAR_53_WIDTH-1:0] ap_iscalar_53_dout,
    output [C_INPUT_SCALAR_54_WIDTH-1:0] ap_iscalar_54_dout,
    output [C_INPUT_SCALAR_55_WIDTH-1:0] ap_iscalar_55_dout,
    output [C_INPUT_SCALAR_56_WIDTH-1:0] ap_iscalar_56_dout,
    output [C_INPUT_SCALAR_57_WIDTH-1:0] ap_iscalar_57_dout,
    output [C_INPUT_SCALAR_58_WIDTH-1:0] ap_iscalar_58_dout,
    output [C_INPUT_SCALAR_59_WIDTH-1:0] ap_iscalar_59_dout,
    output [C_INPUT_SCALAR_60_WIDTH-1:0] ap_iscalar_60_dout,
    output [C_INPUT_SCALAR_61_WIDTH-1:0] ap_iscalar_61_dout,
    output [C_INPUT_SCALAR_62_WIDTH-1:0] ap_iscalar_62_dout,
    output [C_INPUT_SCALAR_63_WIDTH-1:0] ap_iscalar_63_dout,
    output [C_INPUT_SCALAR_64_WIDTH-1:0] ap_iscalar_64_dout,
    output [C_INPUT_SCALAR_65_WIDTH-1:0] ap_iscalar_65_dout,
    output [C_INPUT_SCALAR_66_WIDTH-1:0] ap_iscalar_66_dout,
    output [C_INPUT_SCALAR_67_WIDTH-1:0] ap_iscalar_67_dout,
    output [C_INPUT_SCALAR_68_WIDTH-1:0] ap_iscalar_68_dout,
    output [C_INPUT_SCALAR_69_WIDTH-1:0] ap_iscalar_69_dout,
    output [C_INPUT_SCALAR_70_WIDTH-1:0] ap_iscalar_70_dout,
    output [C_INPUT_SCALAR_71_WIDTH-1:0] ap_iscalar_71_dout,
    output [C_INPUT_SCALAR_72_WIDTH-1:0] ap_iscalar_72_dout,
    output [C_INPUT_SCALAR_73_WIDTH-1:0] ap_iscalar_73_dout,
    output [C_INPUT_SCALAR_74_WIDTH-1:0] ap_iscalar_74_dout,
    output [C_INPUT_SCALAR_75_WIDTH-1:0] ap_iscalar_75_dout,
    output [C_INPUT_SCALAR_76_WIDTH-1:0] ap_iscalar_76_dout,
    output [C_INPUT_SCALAR_77_WIDTH-1:0] ap_iscalar_77_dout,
    output [C_INPUT_SCALAR_78_WIDTH-1:0] ap_iscalar_78_dout,
    output [C_INPUT_SCALAR_79_WIDTH-1:0] ap_iscalar_79_dout,
    output [C_INPUT_SCALAR_80_WIDTH-1:0] ap_iscalar_80_dout,
    output [C_INPUT_SCALAR_81_WIDTH-1:0] ap_iscalar_81_dout,
    output [C_INPUT_SCALAR_82_WIDTH-1:0] ap_iscalar_82_dout,
    output [C_INPUT_SCALAR_83_WIDTH-1:0] ap_iscalar_83_dout,
    output [C_INPUT_SCALAR_84_WIDTH-1:0] ap_iscalar_84_dout,
    output [C_INPUT_SCALAR_85_WIDTH-1:0] ap_iscalar_85_dout,
    output [C_INPUT_SCALAR_86_WIDTH-1:0] ap_iscalar_86_dout,
    output [C_INPUT_SCALAR_87_WIDTH-1:0] ap_iscalar_87_dout,
    output [C_INPUT_SCALAR_88_WIDTH-1:0] ap_iscalar_88_dout,
    output [C_INPUT_SCALAR_89_WIDTH-1:0] ap_iscalar_89_dout,
    output [C_INPUT_SCALAR_90_WIDTH-1:0] ap_iscalar_90_dout,
    output [C_INPUT_SCALAR_91_WIDTH-1:0] ap_iscalar_91_dout,
    output [C_INPUT_SCALAR_92_WIDTH-1:0] ap_iscalar_92_dout,
    output [C_INPUT_SCALAR_93_WIDTH-1:0] ap_iscalar_93_dout,
    output [C_INPUT_SCALAR_94_WIDTH-1:0] ap_iscalar_94_dout,
    output [C_INPUT_SCALAR_95_WIDTH-1:0] ap_iscalar_95_dout,
    output [C_INPUT_SCALAR_96_WIDTH-1:0] ap_iscalar_96_dout,
    output [C_INPUT_SCALAR_97_WIDTH-1:0] ap_iscalar_97_dout,
    output [C_INPUT_SCALAR_98_WIDTH-1:0] ap_iscalar_98_dout,
    output [C_INPUT_SCALAR_99_WIDTH-1:0] ap_iscalar_99_dout,
    output [C_INPUT_SCALAR_100_WIDTH-1:0] ap_iscalar_100_dout,
    output [C_INPUT_SCALAR_101_WIDTH-1:0] ap_iscalar_101_dout,
    output [C_INPUT_SCALAR_102_WIDTH-1:0] ap_iscalar_102_dout,
    output [C_INPUT_SCALAR_103_WIDTH-1:0] ap_iscalar_103_dout,
    output [C_INPUT_SCALAR_104_WIDTH-1:0] ap_iscalar_104_dout,
    output [C_INPUT_SCALAR_105_WIDTH-1:0] ap_iscalar_105_dout,
    output [C_INPUT_SCALAR_106_WIDTH-1:0] ap_iscalar_106_dout,
    output [C_INPUT_SCALAR_107_WIDTH-1:0] ap_iscalar_107_dout,
    output [C_INPUT_SCALAR_108_WIDTH-1:0] ap_iscalar_108_dout,
    output [C_INPUT_SCALAR_109_WIDTH-1:0] ap_iscalar_109_dout,
    output [C_INPUT_SCALAR_110_WIDTH-1:0] ap_iscalar_110_dout,
    output [C_INPUT_SCALAR_111_WIDTH-1:0] ap_iscalar_111_dout,
    output [C_INPUT_SCALAR_112_WIDTH-1:0] ap_iscalar_112_dout,
    output [C_INPUT_SCALAR_113_WIDTH-1:0] ap_iscalar_113_dout,
    output [C_INPUT_SCALAR_114_WIDTH-1:0] ap_iscalar_114_dout,
    output [C_INPUT_SCALAR_115_WIDTH-1:0] ap_iscalar_115_dout,
    output [C_INPUT_SCALAR_116_WIDTH-1:0] ap_iscalar_116_dout,
    output [C_INPUT_SCALAR_117_WIDTH-1:0] ap_iscalar_117_dout,
    output [C_INPUT_SCALAR_118_WIDTH-1:0] ap_iscalar_118_dout,
    output [C_INPUT_SCALAR_119_WIDTH-1:0] ap_iscalar_119_dout,
    output [C_INPUT_SCALAR_120_WIDTH-1:0] ap_iscalar_120_dout,
    output [C_INPUT_SCALAR_121_WIDTH-1:0] ap_iscalar_121_dout,
    output [C_INPUT_SCALAR_122_WIDTH-1:0] ap_iscalar_122_dout,
    output [C_INPUT_SCALAR_123_WIDTH-1:0] ap_iscalar_123_dout,
    output [C_INPUT_SCALAR_124_WIDTH-1:0] ap_iscalar_124_dout,
    output [C_INPUT_SCALAR_125_WIDTH-1:0] ap_iscalar_125_dout,
    output [C_INPUT_SCALAR_126_WIDTH-1:0] ap_iscalar_126_dout,
    output [C_INPUT_SCALAR_127_WIDTH-1:0] ap_iscalar_127_dout,
    //output scalar ports
    input [C_OUTPUT_SCALAR_0_WIDTH-1:0] ap_oscalar_0_din,
    input [C_OUTPUT_SCALAR_1_WIDTH-1:0] ap_oscalar_1_din,
    input [C_OUTPUT_SCALAR_2_WIDTH-1:0] ap_oscalar_2_din,
    input [C_OUTPUT_SCALAR_3_WIDTH-1:0] ap_oscalar_3_din,
    input [C_OUTPUT_SCALAR_4_WIDTH-1:0] ap_oscalar_4_din,
    input [C_OUTPUT_SCALAR_5_WIDTH-1:0] ap_oscalar_5_din,
    input [C_OUTPUT_SCALAR_6_WIDTH-1:0] ap_oscalar_6_din,
    input [C_OUTPUT_SCALAR_7_WIDTH-1:0] ap_oscalar_7_din,
    input [C_OUTPUT_SCALAR_8_WIDTH-1:0] ap_oscalar_8_din,
    input [C_OUTPUT_SCALAR_9_WIDTH-1:0] ap_oscalar_9_din,
    input [C_OUTPUT_SCALAR_10_WIDTH-1:0] ap_oscalar_10_din,
    input [C_OUTPUT_SCALAR_11_WIDTH-1:0] ap_oscalar_11_din,
    input [C_OUTPUT_SCALAR_12_WIDTH-1:0] ap_oscalar_12_din,
    input [C_OUTPUT_SCALAR_13_WIDTH-1:0] ap_oscalar_13_din,
    input [C_OUTPUT_SCALAR_14_WIDTH-1:0] ap_oscalar_14_din,
    input [C_OUTPUT_SCALAR_15_WIDTH-1:0] ap_oscalar_15_din,
    input [C_OUTPUT_SCALAR_16_WIDTH-1:0] ap_oscalar_16_din,
    input [C_OUTPUT_SCALAR_17_WIDTH-1:0] ap_oscalar_17_din,
    input [C_OUTPUT_SCALAR_18_WIDTH-1:0] ap_oscalar_18_din,
    input [C_OUTPUT_SCALAR_19_WIDTH-1:0] ap_oscalar_19_din,
    input [C_OUTPUT_SCALAR_20_WIDTH-1:0] ap_oscalar_20_din,
    input [C_OUTPUT_SCALAR_21_WIDTH-1:0] ap_oscalar_21_din,
    input [C_OUTPUT_SCALAR_22_WIDTH-1:0] ap_oscalar_22_din,
    input [C_OUTPUT_SCALAR_23_WIDTH-1:0] ap_oscalar_23_din,
    input [C_OUTPUT_SCALAR_24_WIDTH-1:0] ap_oscalar_24_din,
    input [C_OUTPUT_SCALAR_25_WIDTH-1:0] ap_oscalar_25_din,
    input [C_OUTPUT_SCALAR_26_WIDTH-1:0] ap_oscalar_26_din,
    input [C_OUTPUT_SCALAR_27_WIDTH-1:0] ap_oscalar_27_din,
    input [C_OUTPUT_SCALAR_28_WIDTH-1:0] ap_oscalar_28_din,
    input [C_OUTPUT_SCALAR_29_WIDTH-1:0] ap_oscalar_29_din,
    input [C_OUTPUT_SCALAR_30_WIDTH-1:0] ap_oscalar_30_din,
    input [C_OUTPUT_SCALAR_31_WIDTH-1:0] ap_oscalar_31_din,
    input [C_OUTPUT_SCALAR_32_WIDTH-1:0] ap_oscalar_32_din,
    input [C_OUTPUT_SCALAR_33_WIDTH-1:0] ap_oscalar_33_din,
    input [C_OUTPUT_SCALAR_34_WIDTH-1:0] ap_oscalar_34_din,
    input [C_OUTPUT_SCALAR_35_WIDTH-1:0] ap_oscalar_35_din,
    input [C_OUTPUT_SCALAR_36_WIDTH-1:0] ap_oscalar_36_din,
    input [C_OUTPUT_SCALAR_37_WIDTH-1:0] ap_oscalar_37_din,
    input [C_OUTPUT_SCALAR_38_WIDTH-1:0] ap_oscalar_38_din,
    input [C_OUTPUT_SCALAR_39_WIDTH-1:0] ap_oscalar_39_din,
    input [C_OUTPUT_SCALAR_40_WIDTH-1:0] ap_oscalar_40_din,
    input [C_OUTPUT_SCALAR_41_WIDTH-1:0] ap_oscalar_41_din,
    input [C_OUTPUT_SCALAR_42_WIDTH-1:0] ap_oscalar_42_din,
    input [C_OUTPUT_SCALAR_43_WIDTH-1:0] ap_oscalar_43_din,
    input [C_OUTPUT_SCALAR_44_WIDTH-1:0] ap_oscalar_44_din,
    input [C_OUTPUT_SCALAR_45_WIDTH-1:0] ap_oscalar_45_din,
    input [C_OUTPUT_SCALAR_46_WIDTH-1:0] ap_oscalar_46_din,
    input [C_OUTPUT_SCALAR_47_WIDTH-1:0] ap_oscalar_47_din,
    input [C_OUTPUT_SCALAR_48_WIDTH-1:0] ap_oscalar_48_din,
    input [C_OUTPUT_SCALAR_49_WIDTH-1:0] ap_oscalar_49_din,
    input [C_OUTPUT_SCALAR_50_WIDTH-1:0] ap_oscalar_50_din,
    input [C_OUTPUT_SCALAR_51_WIDTH-1:0] ap_oscalar_51_din,
    input [C_OUTPUT_SCALAR_52_WIDTH-1:0] ap_oscalar_52_din,
    input [C_OUTPUT_SCALAR_53_WIDTH-1:0] ap_oscalar_53_din,
    input [C_OUTPUT_SCALAR_54_WIDTH-1:0] ap_oscalar_54_din,
    input [C_OUTPUT_SCALAR_55_WIDTH-1:0] ap_oscalar_55_din,
    input [C_OUTPUT_SCALAR_56_WIDTH-1:0] ap_oscalar_56_din,
    input [C_OUTPUT_SCALAR_57_WIDTH-1:0] ap_oscalar_57_din,
    input [C_OUTPUT_SCALAR_58_WIDTH-1:0] ap_oscalar_58_din,
    input [C_OUTPUT_SCALAR_59_WIDTH-1:0] ap_oscalar_59_din,
    input [C_OUTPUT_SCALAR_60_WIDTH-1:0] ap_oscalar_60_din,
    input [C_OUTPUT_SCALAR_61_WIDTH-1:0] ap_oscalar_61_din,
    input [C_OUTPUT_SCALAR_62_WIDTH-1:0] ap_oscalar_62_din,
    input [C_OUTPUT_SCALAR_63_WIDTH-1:0] ap_oscalar_63_din,
    input [C_OUTPUT_SCALAR_64_WIDTH-1:0] ap_oscalar_64_din,
    input [C_OUTPUT_SCALAR_65_WIDTH-1:0] ap_oscalar_65_din,
    input [C_OUTPUT_SCALAR_66_WIDTH-1:0] ap_oscalar_66_din,
    input [C_OUTPUT_SCALAR_67_WIDTH-1:0] ap_oscalar_67_din,
    input [C_OUTPUT_SCALAR_68_WIDTH-1:0] ap_oscalar_68_din,
    input [C_OUTPUT_SCALAR_69_WIDTH-1:0] ap_oscalar_69_din,
    input [C_OUTPUT_SCALAR_70_WIDTH-1:0] ap_oscalar_70_din,
    input [C_OUTPUT_SCALAR_71_WIDTH-1:0] ap_oscalar_71_din,
    input [C_OUTPUT_SCALAR_72_WIDTH-1:0] ap_oscalar_72_din,
    input [C_OUTPUT_SCALAR_73_WIDTH-1:0] ap_oscalar_73_din,
    input [C_OUTPUT_SCALAR_74_WIDTH-1:0] ap_oscalar_74_din,
    input [C_OUTPUT_SCALAR_75_WIDTH-1:0] ap_oscalar_75_din,
    input [C_OUTPUT_SCALAR_76_WIDTH-1:0] ap_oscalar_76_din,
    input [C_OUTPUT_SCALAR_77_WIDTH-1:0] ap_oscalar_77_din,
    input [C_OUTPUT_SCALAR_78_WIDTH-1:0] ap_oscalar_78_din,
    input [C_OUTPUT_SCALAR_79_WIDTH-1:0] ap_oscalar_79_din,
    input [C_OUTPUT_SCALAR_80_WIDTH-1:0] ap_oscalar_80_din,
    input [C_OUTPUT_SCALAR_81_WIDTH-1:0] ap_oscalar_81_din,
    input [C_OUTPUT_SCALAR_82_WIDTH-1:0] ap_oscalar_82_din,
    input [C_OUTPUT_SCALAR_83_WIDTH-1:0] ap_oscalar_83_din,
    input [C_OUTPUT_SCALAR_84_WIDTH-1:0] ap_oscalar_84_din,
    input [C_OUTPUT_SCALAR_85_WIDTH-1:0] ap_oscalar_85_din,
    input [C_OUTPUT_SCALAR_86_WIDTH-1:0] ap_oscalar_86_din,
    input [C_OUTPUT_SCALAR_87_WIDTH-1:0] ap_oscalar_87_din,
    input [C_OUTPUT_SCALAR_88_WIDTH-1:0] ap_oscalar_88_din,
    input [C_OUTPUT_SCALAR_89_WIDTH-1:0] ap_oscalar_89_din,
    input [C_OUTPUT_SCALAR_90_WIDTH-1:0] ap_oscalar_90_din,
    input [C_OUTPUT_SCALAR_91_WIDTH-1:0] ap_oscalar_91_din,
    input [C_OUTPUT_SCALAR_92_WIDTH-1:0] ap_oscalar_92_din,
    input [C_OUTPUT_SCALAR_93_WIDTH-1:0] ap_oscalar_93_din,
    input [C_OUTPUT_SCALAR_94_WIDTH-1:0] ap_oscalar_94_din,
    input [C_OUTPUT_SCALAR_95_WIDTH-1:0] ap_oscalar_95_din,
    input [C_OUTPUT_SCALAR_96_WIDTH-1:0] ap_oscalar_96_din,
    input [C_OUTPUT_SCALAR_97_WIDTH-1:0] ap_oscalar_97_din,
    input [C_OUTPUT_SCALAR_98_WIDTH-1:0] ap_oscalar_98_din,
    input [C_OUTPUT_SCALAR_99_WIDTH-1:0] ap_oscalar_99_din,
    input [C_OUTPUT_SCALAR_100_WIDTH-1:0] ap_oscalar_100_din,
    input [C_OUTPUT_SCALAR_101_WIDTH-1:0] ap_oscalar_101_din,
    input [C_OUTPUT_SCALAR_102_WIDTH-1:0] ap_oscalar_102_din,
    input [C_OUTPUT_SCALAR_103_WIDTH-1:0] ap_oscalar_103_din,
    input [C_OUTPUT_SCALAR_104_WIDTH-1:0] ap_oscalar_104_din,
    input [C_OUTPUT_SCALAR_105_WIDTH-1:0] ap_oscalar_105_din,
    input [C_OUTPUT_SCALAR_106_WIDTH-1:0] ap_oscalar_106_din,
    input [C_OUTPUT_SCALAR_107_WIDTH-1:0] ap_oscalar_107_din,
    input [C_OUTPUT_SCALAR_108_WIDTH-1:0] ap_oscalar_108_din,
    input [C_OUTPUT_SCALAR_109_WIDTH-1:0] ap_oscalar_109_din,
    input [C_OUTPUT_SCALAR_110_WIDTH-1:0] ap_oscalar_110_din,
    input [C_OUTPUT_SCALAR_111_WIDTH-1:0] ap_oscalar_111_din,
    input [C_OUTPUT_SCALAR_112_WIDTH-1:0] ap_oscalar_112_din,
    input [C_OUTPUT_SCALAR_113_WIDTH-1:0] ap_oscalar_113_din,
    input [C_OUTPUT_SCALAR_114_WIDTH-1:0] ap_oscalar_114_din,
    input [C_OUTPUT_SCALAR_115_WIDTH-1:0] ap_oscalar_115_din,
    input [C_OUTPUT_SCALAR_116_WIDTH-1:0] ap_oscalar_116_din,
    input [C_OUTPUT_SCALAR_117_WIDTH-1:0] ap_oscalar_117_din,
    input [C_OUTPUT_SCALAR_118_WIDTH-1:0] ap_oscalar_118_din,
    input [C_OUTPUT_SCALAR_119_WIDTH-1:0] ap_oscalar_119_din,
    input [C_OUTPUT_SCALAR_120_WIDTH-1:0] ap_oscalar_120_din,
    input [C_OUTPUT_SCALAR_121_WIDTH-1:0] ap_oscalar_121_din,
    input [C_OUTPUT_SCALAR_122_WIDTH-1:0] ap_oscalar_122_din,
    input [C_OUTPUT_SCALAR_123_WIDTH-1:0] ap_oscalar_123_din,
    input [C_OUTPUT_SCALAR_124_WIDTH-1:0] ap_oscalar_124_din,
    input [C_OUTPUT_SCALAR_125_WIDTH-1:0] ap_oscalar_125_din,
    input [C_OUTPUT_SCALAR_126_WIDTH-1:0] ap_oscalar_126_din,
    input [C_OUTPUT_SCALAR_127_WIDTH-1:0] ap_oscalar_127_din,
    //output scalar valid ports
    input ap_oscalar_0_vld,
    input ap_oscalar_1_vld,
    input ap_oscalar_2_vld,
    input ap_oscalar_3_vld,
    input ap_oscalar_4_vld,
    input ap_oscalar_5_vld,
    input ap_oscalar_6_vld,
    input ap_oscalar_7_vld,
    input ap_oscalar_8_vld,
    input ap_oscalar_9_vld,
    input ap_oscalar_10_vld,
    input ap_oscalar_11_vld,
    input ap_oscalar_12_vld,
    input ap_oscalar_13_vld,
    input ap_oscalar_14_vld,
    input ap_oscalar_15_vld,
    input ap_oscalar_16_vld,
    input ap_oscalar_17_vld,
    input ap_oscalar_18_vld,
    input ap_oscalar_19_vld,
    input ap_oscalar_20_vld,
    input ap_oscalar_21_vld,
    input ap_oscalar_22_vld,
    input ap_oscalar_23_vld,
    input ap_oscalar_24_vld,
    input ap_oscalar_25_vld,
    input ap_oscalar_26_vld,
    input ap_oscalar_27_vld,
    input ap_oscalar_28_vld,
    input ap_oscalar_29_vld,
    input ap_oscalar_30_vld,
    input ap_oscalar_31_vld,
    input ap_oscalar_32_vld,
    input ap_oscalar_33_vld,
    input ap_oscalar_34_vld,
    input ap_oscalar_35_vld,
    input ap_oscalar_36_vld,
    input ap_oscalar_37_vld,
    input ap_oscalar_38_vld,
    input ap_oscalar_39_vld,
    input ap_oscalar_40_vld,
    input ap_oscalar_41_vld,
    input ap_oscalar_42_vld,
    input ap_oscalar_43_vld,
    input ap_oscalar_44_vld,
    input ap_oscalar_45_vld,
    input ap_oscalar_46_vld,
    input ap_oscalar_47_vld,
    input ap_oscalar_48_vld,
    input ap_oscalar_49_vld,
    input ap_oscalar_50_vld,
    input ap_oscalar_51_vld,
    input ap_oscalar_52_vld,
    input ap_oscalar_53_vld,
    input ap_oscalar_54_vld,
    input ap_oscalar_55_vld,
    input ap_oscalar_56_vld,
    input ap_oscalar_57_vld,
    input ap_oscalar_58_vld,
    input ap_oscalar_59_vld,
    input ap_oscalar_60_vld,
    input ap_oscalar_61_vld,
    input ap_oscalar_62_vld,
    input ap_oscalar_63_vld,
    input ap_oscalar_64_vld,
    input ap_oscalar_65_vld,
    input ap_oscalar_66_vld,
    input ap_oscalar_67_vld,
    input ap_oscalar_68_vld,
    input ap_oscalar_69_vld,
    input ap_oscalar_70_vld,
    input ap_oscalar_71_vld,
    input ap_oscalar_72_vld,
    input ap_oscalar_73_vld,
    input ap_oscalar_74_vld,
    input ap_oscalar_75_vld,
    input ap_oscalar_76_vld,
    input ap_oscalar_77_vld,
    input ap_oscalar_78_vld,
    input ap_oscalar_79_vld,
    input ap_oscalar_80_vld,
    input ap_oscalar_81_vld,
    input ap_oscalar_82_vld,
    input ap_oscalar_83_vld,
    input ap_oscalar_84_vld,
    input ap_oscalar_85_vld,
    input ap_oscalar_86_vld,
    input ap_oscalar_87_vld,
    input ap_oscalar_88_vld,
    input ap_oscalar_89_vld,
    input ap_oscalar_90_vld,
    input ap_oscalar_91_vld,
    input ap_oscalar_92_vld,
    input ap_oscalar_93_vld,
    input ap_oscalar_94_vld,
    input ap_oscalar_95_vld,
    input ap_oscalar_96_vld,
    input ap_oscalar_97_vld,
    input ap_oscalar_98_vld,
    input ap_oscalar_99_vld,
    input ap_oscalar_100_vld,
    input ap_oscalar_101_vld,
    input ap_oscalar_102_vld,
    input ap_oscalar_103_vld,
    input ap_oscalar_104_vld,
    input ap_oscalar_105_vld,
    input ap_oscalar_106_vld,
    input ap_oscalar_107_vld,
    input ap_oscalar_108_vld,
    input ap_oscalar_109_vld,
    input ap_oscalar_110_vld,
    input ap_oscalar_111_vld,
    input ap_oscalar_112_vld,
    input ap_oscalar_113_vld,
    input ap_oscalar_114_vld,
    input ap_oscalar_115_vld,
    input ap_oscalar_116_vld,
    input ap_oscalar_117_vld,
    input ap_oscalar_118_vld,
    input ap_oscalar_119_vld,
    input ap_oscalar_120_vld,
    input ap_oscalar_121_vld,
    input ap_oscalar_122_vld,
    input ap_oscalar_123_vld,
    input ap_oscalar_124_vld,
    input ap_oscalar_125_vld,
    input ap_oscalar_126_vld,
    input ap_oscalar_127_vld,
    //-----------------------------------------------------
    //input AXI-Stream to FIFO interface 0
    input s_axis_fifo_0_tlast,
    input s_axis_fifo_0_tvalid,
    input [C_INPUT_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tkeep,
    input [C_INPUT_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tstrb,
    input [C_INPUT_FIFO_0_DMWIDTH-1:0] s_axis_fifo_0_tdata,
    output s_axis_fifo_0_tready,
    output ap_fifo_iarg_0_empty_n,
    output [C_INPUT_FIFO_0_WIDTH-1:0] ap_fifo_iarg_0_dout,
    input ap_fifo_iarg_0_read,
    //input AXI-Stream to FIFO interface 1
    input s_axis_fifo_1_tlast,
    input s_axis_fifo_1_tvalid,
    input [C_INPUT_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tkeep,
    input [C_INPUT_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tstrb,
    input [C_INPUT_FIFO_1_DMWIDTH-1:0] s_axis_fifo_1_tdata,
    output s_axis_fifo_1_tready,
    output ap_fifo_iarg_1_empty_n,
    output [C_INPUT_FIFO_1_WIDTH-1:0] ap_fifo_iarg_1_dout,
    input ap_fifo_iarg_1_read,
    //input AXI-Stream to FIFO interface 2
    input s_axis_fifo_2_tlast,
    input s_axis_fifo_2_tvalid,
    input [C_INPUT_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tkeep,
    input [C_INPUT_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tstrb,
    input [C_INPUT_FIFO_2_DMWIDTH-1:0] s_axis_fifo_2_tdata,
    output s_axis_fifo_2_tready,
    output ap_fifo_iarg_2_empty_n,
    output [C_INPUT_FIFO_2_WIDTH-1:0] ap_fifo_iarg_2_dout,
    input ap_fifo_iarg_2_read,
    //input AXI-Stream to FIFO interface 3
    input s_axis_fifo_3_tlast,
    input s_axis_fifo_3_tvalid,
    input [C_INPUT_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tkeep,
    input [C_INPUT_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tstrb,
    input [C_INPUT_FIFO_3_DMWIDTH-1:0] s_axis_fifo_3_tdata,
    output s_axis_fifo_3_tready,
    output ap_fifo_iarg_3_empty_n,
    output [C_INPUT_FIFO_3_WIDTH-1:0] ap_fifo_iarg_3_dout,
    input ap_fifo_iarg_3_read,
    //input AXI-Stream to FIFO interface 4
    input s_axis_fifo_4_tlast,
    input s_axis_fifo_4_tvalid,
    input [C_INPUT_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tkeep,
    input [C_INPUT_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tstrb,
    input [C_INPUT_FIFO_4_DMWIDTH-1:0] s_axis_fifo_4_tdata,
    output s_axis_fifo_4_tready,
    output ap_fifo_iarg_4_empty_n,
    output [C_INPUT_FIFO_4_WIDTH-1:0] ap_fifo_iarg_4_dout,
    input ap_fifo_iarg_4_read,
    //input AXI-Stream to FIFO interface 5
    input s_axis_fifo_5_tlast,
    input s_axis_fifo_5_tvalid,
    input [C_INPUT_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tkeep,
    input [C_INPUT_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tstrb,
    input [C_INPUT_FIFO_5_DMWIDTH-1:0] s_axis_fifo_5_tdata,
    output s_axis_fifo_5_tready,
    output ap_fifo_iarg_5_empty_n,
    output [C_INPUT_FIFO_5_WIDTH-1:0] ap_fifo_iarg_5_dout,
    input ap_fifo_iarg_5_read,
    //input AXI-Stream to FIFO interface 6
    input s_axis_fifo_6_tlast,
    input s_axis_fifo_6_tvalid,
    input [C_INPUT_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tkeep,
    input [C_INPUT_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tstrb,
    input [C_INPUT_FIFO_6_DMWIDTH-1:0] s_axis_fifo_6_tdata,
    output s_axis_fifo_6_tready,
    output ap_fifo_iarg_6_empty_n,
    output [C_INPUT_FIFO_6_WIDTH-1:0] ap_fifo_iarg_6_dout,
    input ap_fifo_iarg_6_read,
    //input AXI-Stream to FIFO interface 7
    input s_axis_fifo_7_tlast,
    input s_axis_fifo_7_tvalid,
    input [C_INPUT_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tkeep,
    input [C_INPUT_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tstrb,
    input [C_INPUT_FIFO_7_DMWIDTH-1:0] s_axis_fifo_7_tdata,
    output s_axis_fifo_7_tready,
    output ap_fifo_iarg_7_empty_n,
    output [C_INPUT_FIFO_7_WIDTH-1:0] ap_fifo_iarg_7_dout,
    input ap_fifo_iarg_7_read,
    //input AXI-Stream to FIFO interface 8
    input s_axis_fifo_8_tlast,
    input s_axis_fifo_8_tvalid,
    input [C_INPUT_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tkeep,
    input [C_INPUT_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tstrb,
    input [C_INPUT_FIFO_8_DMWIDTH-1:0] s_axis_fifo_8_tdata,
    output s_axis_fifo_8_tready,
    output ap_fifo_iarg_8_empty_n,
    output [C_INPUT_FIFO_8_WIDTH-1:0] ap_fifo_iarg_8_dout,
    input ap_fifo_iarg_8_read,
    //input AXI-Stream to FIFO interface 9
    input s_axis_fifo_9_tlast,
    input s_axis_fifo_9_tvalid,
    input [C_INPUT_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tkeep,
    input [C_INPUT_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tstrb,
    input [C_INPUT_FIFO_9_DMWIDTH-1:0] s_axis_fifo_9_tdata,
    output s_axis_fifo_9_tready,
    output ap_fifo_iarg_9_empty_n,
    output [C_INPUT_FIFO_9_WIDTH-1:0] ap_fifo_iarg_9_dout,
    input ap_fifo_iarg_9_read,
    //input AXI-Stream to FIFO interface 10
    input s_axis_fifo_10_tlast,
    input s_axis_fifo_10_tvalid,
    input [C_INPUT_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tkeep,
    input [C_INPUT_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tstrb,
    input [C_INPUT_FIFO_10_DMWIDTH-1:0] s_axis_fifo_10_tdata,
    output s_axis_fifo_10_tready,
    output ap_fifo_iarg_10_empty_n,
    output [C_INPUT_FIFO_10_WIDTH-1:0] ap_fifo_iarg_10_dout,
    input ap_fifo_iarg_10_read,
    //input AXI-Stream to FIFO interface 11
    input s_axis_fifo_11_tlast,
    input s_axis_fifo_11_tvalid,
    input [C_INPUT_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tkeep,
    input [C_INPUT_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tstrb,
    input [C_INPUT_FIFO_11_DMWIDTH-1:0] s_axis_fifo_11_tdata,
    output s_axis_fifo_11_tready,
    output ap_fifo_iarg_11_empty_n,
    output [C_INPUT_FIFO_11_WIDTH-1:0] ap_fifo_iarg_11_dout,
    input ap_fifo_iarg_11_read,
    //input AXI-Stream to FIFO interface 12
    input s_axis_fifo_12_tlast,
    input s_axis_fifo_12_tvalid,
    input [C_INPUT_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tkeep,
    input [C_INPUT_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tstrb,
    input [C_INPUT_FIFO_12_DMWIDTH-1:0] s_axis_fifo_12_tdata,
    output s_axis_fifo_12_tready,
    output ap_fifo_iarg_12_empty_n,
    output [C_INPUT_FIFO_12_WIDTH-1:0] ap_fifo_iarg_12_dout,
    input ap_fifo_iarg_12_read,
    //input AXI-Stream to FIFO interface 13
    input s_axis_fifo_13_tlast,
    input s_axis_fifo_13_tvalid,
    input [C_INPUT_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tkeep,
    input [C_INPUT_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tstrb,
    input [C_INPUT_FIFO_13_DMWIDTH-1:0] s_axis_fifo_13_tdata,
    output s_axis_fifo_13_tready,
    output ap_fifo_iarg_13_empty_n,
    output [C_INPUT_FIFO_13_WIDTH-1:0] ap_fifo_iarg_13_dout,
    input ap_fifo_iarg_13_read,
    //input AXI-Stream to FIFO interface 14
    input s_axis_fifo_14_tlast,
    input s_axis_fifo_14_tvalid,
    input [C_INPUT_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tkeep,
    input [C_INPUT_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tstrb,
    input [C_INPUT_FIFO_14_DMWIDTH-1:0] s_axis_fifo_14_tdata,
    output s_axis_fifo_14_tready,
    output ap_fifo_iarg_14_empty_n,
    output [C_INPUT_FIFO_14_WIDTH-1:0] ap_fifo_iarg_14_dout,
    input ap_fifo_iarg_14_read,
    //input AXI-Stream to FIFO interface 15
    input s_axis_fifo_15_tlast,
    input s_axis_fifo_15_tvalid,
    input [C_INPUT_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tkeep,
    input [C_INPUT_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tstrb,
    input [C_INPUT_FIFO_15_DMWIDTH-1:0] s_axis_fifo_15_tdata,
    output s_axis_fifo_15_tready,
    output ap_fifo_iarg_15_empty_n,
    output [C_INPUT_FIFO_15_WIDTH-1:0] ap_fifo_iarg_15_dout,
    input ap_fifo_iarg_15_read,
    //input AXI-Stream to FIFO interface 16
    input s_axis_fifo_16_tlast,
    input s_axis_fifo_16_tvalid,
    input [C_INPUT_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tkeep,
    input [C_INPUT_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tstrb,
    input [C_INPUT_FIFO_16_DMWIDTH-1:0] s_axis_fifo_16_tdata,
    output s_axis_fifo_16_tready,
    output ap_fifo_iarg_16_empty_n,
    output [C_INPUT_FIFO_16_WIDTH-1:0] ap_fifo_iarg_16_dout,
    input ap_fifo_iarg_16_read,
    //input AXI-Stream to FIFO interface 17
    input s_axis_fifo_17_tlast,
    input s_axis_fifo_17_tvalid,
    input [C_INPUT_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tkeep,
    input [C_INPUT_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tstrb,
    input [C_INPUT_FIFO_17_DMWIDTH-1:0] s_axis_fifo_17_tdata,
    output s_axis_fifo_17_tready,
    output ap_fifo_iarg_17_empty_n,
    output [C_INPUT_FIFO_17_WIDTH-1:0] ap_fifo_iarg_17_dout,
    input ap_fifo_iarg_17_read,
    //input AXI-Stream to FIFO interface 18
    input s_axis_fifo_18_tlast,
    input s_axis_fifo_18_tvalid,
    input [C_INPUT_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tkeep,
    input [C_INPUT_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tstrb,
    input [C_INPUT_FIFO_18_DMWIDTH-1:0] s_axis_fifo_18_tdata,
    output s_axis_fifo_18_tready,
    output ap_fifo_iarg_18_empty_n,
    output [C_INPUT_FIFO_18_WIDTH-1:0] ap_fifo_iarg_18_dout,
    input ap_fifo_iarg_18_read,
    //input AXI-Stream to FIFO interface 19
    input s_axis_fifo_19_tlast,
    input s_axis_fifo_19_tvalid,
    input [C_INPUT_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tkeep,
    input [C_INPUT_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tstrb,
    input [C_INPUT_FIFO_19_DMWIDTH-1:0] s_axis_fifo_19_tdata,
    output s_axis_fifo_19_tready,
    output ap_fifo_iarg_19_empty_n,
    output [C_INPUT_FIFO_19_WIDTH-1:0] ap_fifo_iarg_19_dout,
    input ap_fifo_iarg_19_read,
    //input AXI-Stream to FIFO interface 20
    input s_axis_fifo_20_tlast,
    input s_axis_fifo_20_tvalid,
    input [C_INPUT_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tkeep,
    input [C_INPUT_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tstrb,
    input [C_INPUT_FIFO_20_DMWIDTH-1:0] s_axis_fifo_20_tdata,
    output s_axis_fifo_20_tready,
    output ap_fifo_iarg_20_empty_n,
    output [C_INPUT_FIFO_20_WIDTH-1:0] ap_fifo_iarg_20_dout,
    input ap_fifo_iarg_20_read,
    //input AXI-Stream to FIFO interface 21
    input s_axis_fifo_21_tlast,
    input s_axis_fifo_21_tvalid,
    input [C_INPUT_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tkeep,
    input [C_INPUT_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tstrb,
    input [C_INPUT_FIFO_21_DMWIDTH-1:0] s_axis_fifo_21_tdata,
    output s_axis_fifo_21_tready,
    output ap_fifo_iarg_21_empty_n,
    output [C_INPUT_FIFO_21_WIDTH-1:0] ap_fifo_iarg_21_dout,
    input ap_fifo_iarg_21_read,
    //input AXI-Stream to FIFO interface 22
    input s_axis_fifo_22_tlast,
    input s_axis_fifo_22_tvalid,
    input [C_INPUT_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tkeep,
    input [C_INPUT_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tstrb,
    input [C_INPUT_FIFO_22_DMWIDTH-1:0] s_axis_fifo_22_tdata,
    output s_axis_fifo_22_tready,
    output ap_fifo_iarg_22_empty_n,
    output [C_INPUT_FIFO_22_WIDTH-1:0] ap_fifo_iarg_22_dout,
    input ap_fifo_iarg_22_read,
    //input AXI-Stream to FIFO interface 23
    input s_axis_fifo_23_tlast,
    input s_axis_fifo_23_tvalid,
    input [C_INPUT_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tkeep,
    input [C_INPUT_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tstrb,
    input [C_INPUT_FIFO_23_DMWIDTH-1:0] s_axis_fifo_23_tdata,
    output s_axis_fifo_23_tready,
    output ap_fifo_iarg_23_empty_n,
    output [C_INPUT_FIFO_23_WIDTH-1:0] ap_fifo_iarg_23_dout,
    input ap_fifo_iarg_23_read,
    //input AXI-Stream to FIFO interface 24
    input s_axis_fifo_24_tlast,
    input s_axis_fifo_24_tvalid,
    input [C_INPUT_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tkeep,
    input [C_INPUT_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tstrb,
    input [C_INPUT_FIFO_24_DMWIDTH-1:0] s_axis_fifo_24_tdata,
    output s_axis_fifo_24_tready,
    output ap_fifo_iarg_24_empty_n,
    output [C_INPUT_FIFO_24_WIDTH-1:0] ap_fifo_iarg_24_dout,
    input ap_fifo_iarg_24_read,
    //input AXI-Stream to FIFO interface 25
    input s_axis_fifo_25_tlast,
    input s_axis_fifo_25_tvalid,
    input [C_INPUT_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tkeep,
    input [C_INPUT_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tstrb,
    input [C_INPUT_FIFO_25_DMWIDTH-1:0] s_axis_fifo_25_tdata,
    output s_axis_fifo_25_tready,
    output ap_fifo_iarg_25_empty_n,
    output [C_INPUT_FIFO_25_WIDTH-1:0] ap_fifo_iarg_25_dout,
    input ap_fifo_iarg_25_read,
    //input AXI-Stream to FIFO interface 26
    input s_axis_fifo_26_tlast,
    input s_axis_fifo_26_tvalid,
    input [C_INPUT_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tkeep,
    input [C_INPUT_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tstrb,
    input [C_INPUT_FIFO_26_DMWIDTH-1:0] s_axis_fifo_26_tdata,
    output s_axis_fifo_26_tready,
    output ap_fifo_iarg_26_empty_n,
    output [C_INPUT_FIFO_26_WIDTH-1:0] ap_fifo_iarg_26_dout,
    input ap_fifo_iarg_26_read,
    //input AXI-Stream to FIFO interface 27
    input s_axis_fifo_27_tlast,
    input s_axis_fifo_27_tvalid,
    input [C_INPUT_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tkeep,
    input [C_INPUT_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tstrb,
    input [C_INPUT_FIFO_27_DMWIDTH-1:0] s_axis_fifo_27_tdata,
    output s_axis_fifo_27_tready,
    output ap_fifo_iarg_27_empty_n,
    output [C_INPUT_FIFO_27_WIDTH-1:0] ap_fifo_iarg_27_dout,
    input ap_fifo_iarg_27_read,
    //input AXI-Stream to FIFO interface 28
    input s_axis_fifo_28_tlast,
    input s_axis_fifo_28_tvalid,
    input [C_INPUT_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tkeep,
    input [C_INPUT_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tstrb,
    input [C_INPUT_FIFO_28_DMWIDTH-1:0] s_axis_fifo_28_tdata,
    output s_axis_fifo_28_tready,
    output ap_fifo_iarg_28_empty_n,
    output [C_INPUT_FIFO_28_WIDTH-1:0] ap_fifo_iarg_28_dout,
    input ap_fifo_iarg_28_read,
    //input AXI-Stream to FIFO interface 29
    input s_axis_fifo_29_tlast,
    input s_axis_fifo_29_tvalid,
    input [C_INPUT_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tkeep,
    input [C_INPUT_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tstrb,
    input [C_INPUT_FIFO_29_DMWIDTH-1:0] s_axis_fifo_29_tdata,
    output s_axis_fifo_29_tready,
    output ap_fifo_iarg_29_empty_n,
    output [C_INPUT_FIFO_29_WIDTH-1:0] ap_fifo_iarg_29_dout,
    input ap_fifo_iarg_29_read,
    //input AXI-Stream to FIFO interface 30
    input s_axis_fifo_30_tlast,
    input s_axis_fifo_30_tvalid,
    input [C_INPUT_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tkeep,
    input [C_INPUT_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tstrb,
    input [C_INPUT_FIFO_30_DMWIDTH-1:0] s_axis_fifo_30_tdata,
    output s_axis_fifo_30_tready,
    output ap_fifo_iarg_30_empty_n,
    output [C_INPUT_FIFO_30_WIDTH-1:0] ap_fifo_iarg_30_dout,
    input ap_fifo_iarg_30_read,
    //input AXI-Stream to FIFO interface 31
    input s_axis_fifo_31_tlast,
    input s_axis_fifo_31_tvalid,
    input [C_INPUT_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tkeep,
    input [C_INPUT_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tstrb,
    input [C_INPUT_FIFO_31_DMWIDTH-1:0] s_axis_fifo_31_tdata,
    output s_axis_fifo_31_tready,
    output ap_fifo_iarg_31_empty_n,
    output [C_INPUT_FIFO_31_WIDTH-1:0] ap_fifo_iarg_31_dout,
    input ap_fifo_iarg_31_read,
    //input AXI-Stream to FIFO interface 32
    input s_axis_fifo_32_tlast,
    input s_axis_fifo_32_tvalid,
    input [C_INPUT_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tkeep,
    input [C_INPUT_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tstrb,
    input [C_INPUT_FIFO_32_DMWIDTH-1:0] s_axis_fifo_32_tdata,
    output s_axis_fifo_32_tready,
    output ap_fifo_iarg_32_empty_n,
    output [C_INPUT_FIFO_32_WIDTH-1:0] ap_fifo_iarg_32_dout,
    input ap_fifo_iarg_32_read,
    //input AXI-Stream to FIFO interface 33
    input s_axis_fifo_33_tlast,
    input s_axis_fifo_33_tvalid,
    input [C_INPUT_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tkeep,
    input [C_INPUT_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tstrb,
    input [C_INPUT_FIFO_33_DMWIDTH-1:0] s_axis_fifo_33_tdata,
    output s_axis_fifo_33_tready,
    output ap_fifo_iarg_33_empty_n,
    output [C_INPUT_FIFO_33_WIDTH-1:0] ap_fifo_iarg_33_dout,
    input ap_fifo_iarg_33_read,
    //input AXI-Stream to FIFO interface 34
    input s_axis_fifo_34_tlast,
    input s_axis_fifo_34_tvalid,
    input [C_INPUT_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tkeep,
    input [C_INPUT_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tstrb,
    input [C_INPUT_FIFO_34_DMWIDTH-1:0] s_axis_fifo_34_tdata,
    output s_axis_fifo_34_tready,
    output ap_fifo_iarg_34_empty_n,
    output [C_INPUT_FIFO_34_WIDTH-1:0] ap_fifo_iarg_34_dout,
    input ap_fifo_iarg_34_read,
    //input AXI-Stream to FIFO interface 35
    input s_axis_fifo_35_tlast,
    input s_axis_fifo_35_tvalid,
    input [C_INPUT_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tkeep,
    input [C_INPUT_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tstrb,
    input [C_INPUT_FIFO_35_DMWIDTH-1:0] s_axis_fifo_35_tdata,
    output s_axis_fifo_35_tready,
    output ap_fifo_iarg_35_empty_n,
    output [C_INPUT_FIFO_35_WIDTH-1:0] ap_fifo_iarg_35_dout,
    input ap_fifo_iarg_35_read,
    //input AXI-Stream to FIFO interface 36
    input s_axis_fifo_36_tlast,
    input s_axis_fifo_36_tvalid,
    input [C_INPUT_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tkeep,
    input [C_INPUT_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tstrb,
    input [C_INPUT_FIFO_36_DMWIDTH-1:0] s_axis_fifo_36_tdata,
    output s_axis_fifo_36_tready,
    output ap_fifo_iarg_36_empty_n,
    output [C_INPUT_FIFO_36_WIDTH-1:0] ap_fifo_iarg_36_dout,
    input ap_fifo_iarg_36_read,
    //input AXI-Stream to FIFO interface 37
    input s_axis_fifo_37_tlast,
    input s_axis_fifo_37_tvalid,
    input [C_INPUT_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tkeep,
    input [C_INPUT_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tstrb,
    input [C_INPUT_FIFO_37_DMWIDTH-1:0] s_axis_fifo_37_tdata,
    output s_axis_fifo_37_tready,
    output ap_fifo_iarg_37_empty_n,
    output [C_INPUT_FIFO_37_WIDTH-1:0] ap_fifo_iarg_37_dout,
    input ap_fifo_iarg_37_read,
    //input AXI-Stream to FIFO interface 38
    input s_axis_fifo_38_tlast,
    input s_axis_fifo_38_tvalid,
    input [C_INPUT_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tkeep,
    input [C_INPUT_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tstrb,
    input [C_INPUT_FIFO_38_DMWIDTH-1:0] s_axis_fifo_38_tdata,
    output s_axis_fifo_38_tready,
    output ap_fifo_iarg_38_empty_n,
    output [C_INPUT_FIFO_38_WIDTH-1:0] ap_fifo_iarg_38_dout,
    input ap_fifo_iarg_38_read,
    //input AXI-Stream to FIFO interface 39
    input s_axis_fifo_39_tlast,
    input s_axis_fifo_39_tvalid,
    input [C_INPUT_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tkeep,
    input [C_INPUT_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tstrb,
    input [C_INPUT_FIFO_39_DMWIDTH-1:0] s_axis_fifo_39_tdata,
    output s_axis_fifo_39_tready,
    output ap_fifo_iarg_39_empty_n,
    output [C_INPUT_FIFO_39_WIDTH-1:0] ap_fifo_iarg_39_dout,
    input ap_fifo_iarg_39_read,
    //input AXI-Stream to FIFO interface 40
    input s_axis_fifo_40_tlast,
    input s_axis_fifo_40_tvalid,
    input [C_INPUT_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tkeep,
    input [C_INPUT_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tstrb,
    input [C_INPUT_FIFO_40_DMWIDTH-1:0] s_axis_fifo_40_tdata,
    output s_axis_fifo_40_tready,
    output ap_fifo_iarg_40_empty_n,
    output [C_INPUT_FIFO_40_WIDTH-1:0] ap_fifo_iarg_40_dout,
    input ap_fifo_iarg_40_read,
    //input AXI-Stream to FIFO interface 41
    input s_axis_fifo_41_tlast,
    input s_axis_fifo_41_tvalid,
    input [C_INPUT_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tkeep,
    input [C_INPUT_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tstrb,
    input [C_INPUT_FIFO_41_DMWIDTH-1:0] s_axis_fifo_41_tdata,
    output s_axis_fifo_41_tready,
    output ap_fifo_iarg_41_empty_n,
    output [C_INPUT_FIFO_41_WIDTH-1:0] ap_fifo_iarg_41_dout,
    input ap_fifo_iarg_41_read,
    //input AXI-Stream to FIFO interface 42
    input s_axis_fifo_42_tlast,
    input s_axis_fifo_42_tvalid,
    input [C_INPUT_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tkeep,
    input [C_INPUT_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tstrb,
    input [C_INPUT_FIFO_42_DMWIDTH-1:0] s_axis_fifo_42_tdata,
    output s_axis_fifo_42_tready,
    output ap_fifo_iarg_42_empty_n,
    output [C_INPUT_FIFO_42_WIDTH-1:0] ap_fifo_iarg_42_dout,
    input ap_fifo_iarg_42_read,
    //input AXI-Stream to FIFO interface 43
    input s_axis_fifo_43_tlast,
    input s_axis_fifo_43_tvalid,
    input [C_INPUT_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tkeep,
    input [C_INPUT_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tstrb,
    input [C_INPUT_FIFO_43_DMWIDTH-1:0] s_axis_fifo_43_tdata,
    output s_axis_fifo_43_tready,
    output ap_fifo_iarg_43_empty_n,
    output [C_INPUT_FIFO_43_WIDTH-1:0] ap_fifo_iarg_43_dout,
    input ap_fifo_iarg_43_read,
    //input AXI-Stream to FIFO interface 44
    input s_axis_fifo_44_tlast,
    input s_axis_fifo_44_tvalid,
    input [C_INPUT_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tkeep,
    input [C_INPUT_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tstrb,
    input [C_INPUT_FIFO_44_DMWIDTH-1:0] s_axis_fifo_44_tdata,
    output s_axis_fifo_44_tready,
    output ap_fifo_iarg_44_empty_n,
    output [C_INPUT_FIFO_44_WIDTH-1:0] ap_fifo_iarg_44_dout,
    input ap_fifo_iarg_44_read,
    //input AXI-Stream to FIFO interface 45
    input s_axis_fifo_45_tlast,
    input s_axis_fifo_45_tvalid,
    input [C_INPUT_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tkeep,
    input [C_INPUT_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tstrb,
    input [C_INPUT_FIFO_45_DMWIDTH-1:0] s_axis_fifo_45_tdata,
    output s_axis_fifo_45_tready,
    output ap_fifo_iarg_45_empty_n,
    output [C_INPUT_FIFO_45_WIDTH-1:0] ap_fifo_iarg_45_dout,
    input ap_fifo_iarg_45_read,
    //input AXI-Stream to FIFO interface 46
    input s_axis_fifo_46_tlast,
    input s_axis_fifo_46_tvalid,
    input [C_INPUT_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tkeep,
    input [C_INPUT_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tstrb,
    input [C_INPUT_FIFO_46_DMWIDTH-1:0] s_axis_fifo_46_tdata,
    output s_axis_fifo_46_tready,
    output ap_fifo_iarg_46_empty_n,
    output [C_INPUT_FIFO_46_WIDTH-1:0] ap_fifo_iarg_46_dout,
    input ap_fifo_iarg_46_read,
    //input AXI-Stream to FIFO interface 47
    input s_axis_fifo_47_tlast,
    input s_axis_fifo_47_tvalid,
    input [C_INPUT_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tkeep,
    input [C_INPUT_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tstrb,
    input [C_INPUT_FIFO_47_DMWIDTH-1:0] s_axis_fifo_47_tdata,
    output s_axis_fifo_47_tready,
    output ap_fifo_iarg_47_empty_n,
    output [C_INPUT_FIFO_47_WIDTH-1:0] ap_fifo_iarg_47_dout,
    input ap_fifo_iarg_47_read,
    //input AXI-Stream to FIFO interface 48
    input s_axis_fifo_48_tlast,
    input s_axis_fifo_48_tvalid,
    input [C_INPUT_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tkeep,
    input [C_INPUT_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tstrb,
    input [C_INPUT_FIFO_48_DMWIDTH-1:0] s_axis_fifo_48_tdata,
    output s_axis_fifo_48_tready,
    output ap_fifo_iarg_48_empty_n,
    output [C_INPUT_FIFO_48_WIDTH-1:0] ap_fifo_iarg_48_dout,
    input ap_fifo_iarg_48_read,
    //input AXI-Stream to FIFO interface 49
    input s_axis_fifo_49_tlast,
    input s_axis_fifo_49_tvalid,
    input [C_INPUT_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tkeep,
    input [C_INPUT_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tstrb,
    input [C_INPUT_FIFO_49_DMWIDTH-1:0] s_axis_fifo_49_tdata,
    output s_axis_fifo_49_tready,
    output ap_fifo_iarg_49_empty_n,
    output [C_INPUT_FIFO_49_WIDTH-1:0] ap_fifo_iarg_49_dout,
    input ap_fifo_iarg_49_read,
    //input AXI-Stream to FIFO interface 50
    input s_axis_fifo_50_tlast,
    input s_axis_fifo_50_tvalid,
    input [C_INPUT_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tkeep,
    input [C_INPUT_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tstrb,
    input [C_INPUT_FIFO_50_DMWIDTH-1:0] s_axis_fifo_50_tdata,
    output s_axis_fifo_50_tready,
    output ap_fifo_iarg_50_empty_n,
    output [C_INPUT_FIFO_50_WIDTH-1:0] ap_fifo_iarg_50_dout,
    input ap_fifo_iarg_50_read,
    //input AXI-Stream to FIFO interface 51
    input s_axis_fifo_51_tlast,
    input s_axis_fifo_51_tvalid,
    input [C_INPUT_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tkeep,
    input [C_INPUT_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tstrb,
    input [C_INPUT_FIFO_51_DMWIDTH-1:0] s_axis_fifo_51_tdata,
    output s_axis_fifo_51_tready,
    output ap_fifo_iarg_51_empty_n,
    output [C_INPUT_FIFO_51_WIDTH-1:0] ap_fifo_iarg_51_dout,
    input ap_fifo_iarg_51_read,
    //input AXI-Stream to FIFO interface 52
    input s_axis_fifo_52_tlast,
    input s_axis_fifo_52_tvalid,
    input [C_INPUT_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tkeep,
    input [C_INPUT_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tstrb,
    input [C_INPUT_FIFO_52_DMWIDTH-1:0] s_axis_fifo_52_tdata,
    output s_axis_fifo_52_tready,
    output ap_fifo_iarg_52_empty_n,
    output [C_INPUT_FIFO_52_WIDTH-1:0] ap_fifo_iarg_52_dout,
    input ap_fifo_iarg_52_read,
    //input AXI-Stream to FIFO interface 53
    input s_axis_fifo_53_tlast,
    input s_axis_fifo_53_tvalid,
    input [C_INPUT_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tkeep,
    input [C_INPUT_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tstrb,
    input [C_INPUT_FIFO_53_DMWIDTH-1:0] s_axis_fifo_53_tdata,
    output s_axis_fifo_53_tready,
    output ap_fifo_iarg_53_empty_n,
    output [C_INPUT_FIFO_53_WIDTH-1:0] ap_fifo_iarg_53_dout,
    input ap_fifo_iarg_53_read,
    //input AXI-Stream to FIFO interface 54
    input s_axis_fifo_54_tlast,
    input s_axis_fifo_54_tvalid,
    input [C_INPUT_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tkeep,
    input [C_INPUT_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tstrb,
    input [C_INPUT_FIFO_54_DMWIDTH-1:0] s_axis_fifo_54_tdata,
    output s_axis_fifo_54_tready,
    output ap_fifo_iarg_54_empty_n,
    output [C_INPUT_FIFO_54_WIDTH-1:0] ap_fifo_iarg_54_dout,
    input ap_fifo_iarg_54_read,
    //input AXI-Stream to FIFO interface 55
    input s_axis_fifo_55_tlast,
    input s_axis_fifo_55_tvalid,
    input [C_INPUT_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tkeep,
    input [C_INPUT_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tstrb,
    input [C_INPUT_FIFO_55_DMWIDTH-1:0] s_axis_fifo_55_tdata,
    output s_axis_fifo_55_tready,
    output ap_fifo_iarg_55_empty_n,
    output [C_INPUT_FIFO_55_WIDTH-1:0] ap_fifo_iarg_55_dout,
    input ap_fifo_iarg_55_read,
    //input AXI-Stream to FIFO interface 56
    input s_axis_fifo_56_tlast,
    input s_axis_fifo_56_tvalid,
    input [C_INPUT_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tkeep,
    input [C_INPUT_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tstrb,
    input [C_INPUT_FIFO_56_DMWIDTH-1:0] s_axis_fifo_56_tdata,
    output s_axis_fifo_56_tready,
    output ap_fifo_iarg_56_empty_n,
    output [C_INPUT_FIFO_56_WIDTH-1:0] ap_fifo_iarg_56_dout,
    input ap_fifo_iarg_56_read,
    //input AXI-Stream to FIFO interface 57
    input s_axis_fifo_57_tlast,
    input s_axis_fifo_57_tvalid,
    input [C_INPUT_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tkeep,
    input [C_INPUT_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tstrb,
    input [C_INPUT_FIFO_57_DMWIDTH-1:0] s_axis_fifo_57_tdata,
    output s_axis_fifo_57_tready,
    output ap_fifo_iarg_57_empty_n,
    output [C_INPUT_FIFO_57_WIDTH-1:0] ap_fifo_iarg_57_dout,
    input ap_fifo_iarg_57_read,
    //input AXI-Stream to FIFO interface 58
    input s_axis_fifo_58_tlast,
    input s_axis_fifo_58_tvalid,
    input [C_INPUT_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tkeep,
    input [C_INPUT_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tstrb,
    input [C_INPUT_FIFO_58_DMWIDTH-1:0] s_axis_fifo_58_tdata,
    output s_axis_fifo_58_tready,
    output ap_fifo_iarg_58_empty_n,
    output [C_INPUT_FIFO_58_WIDTH-1:0] ap_fifo_iarg_58_dout,
    input ap_fifo_iarg_58_read,
    //input AXI-Stream to FIFO interface 59
    input s_axis_fifo_59_tlast,
    input s_axis_fifo_59_tvalid,
    input [C_INPUT_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tkeep,
    input [C_INPUT_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tstrb,
    input [C_INPUT_FIFO_59_DMWIDTH-1:0] s_axis_fifo_59_tdata,
    output s_axis_fifo_59_tready,
    output ap_fifo_iarg_59_empty_n,
    output [C_INPUT_FIFO_59_WIDTH-1:0] ap_fifo_iarg_59_dout,
    input ap_fifo_iarg_59_read,
    //input AXI-Stream to FIFO interface 60
    input s_axis_fifo_60_tlast,
    input s_axis_fifo_60_tvalid,
    input [C_INPUT_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tkeep,
    input [C_INPUT_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tstrb,
    input [C_INPUT_FIFO_60_DMWIDTH-1:0] s_axis_fifo_60_tdata,
    output s_axis_fifo_60_tready,
    output ap_fifo_iarg_60_empty_n,
    output [C_INPUT_FIFO_60_WIDTH-1:0] ap_fifo_iarg_60_dout,
    input ap_fifo_iarg_60_read,
    //input AXI-Stream to FIFO interface 61
    input s_axis_fifo_61_tlast,
    input s_axis_fifo_61_tvalid,
    input [C_INPUT_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tkeep,
    input [C_INPUT_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tstrb,
    input [C_INPUT_FIFO_61_DMWIDTH-1:0] s_axis_fifo_61_tdata,
    output s_axis_fifo_61_tready,
    output ap_fifo_iarg_61_empty_n,
    output [C_INPUT_FIFO_61_WIDTH-1:0] ap_fifo_iarg_61_dout,
    input ap_fifo_iarg_61_read,
    //input AXI-Stream to FIFO interface 62
    input s_axis_fifo_62_tlast,
    input s_axis_fifo_62_tvalid,
    input [C_INPUT_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tkeep,
    input [C_INPUT_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tstrb,
    input [C_INPUT_FIFO_62_DMWIDTH-1:0] s_axis_fifo_62_tdata,
    output s_axis_fifo_62_tready,
    output ap_fifo_iarg_62_empty_n,
    output [C_INPUT_FIFO_62_WIDTH-1:0] ap_fifo_iarg_62_dout,
    input ap_fifo_iarg_62_read,
    //input AXI-Stream to FIFO interface 63
    input s_axis_fifo_63_tlast,
    input s_axis_fifo_63_tvalid,
    input [C_INPUT_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tkeep,
    input [C_INPUT_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tstrb,
    input [C_INPUT_FIFO_63_DMWIDTH-1:0] s_axis_fifo_63_tdata,
    output s_axis_fifo_63_tready,
    output ap_fifo_iarg_63_empty_n,
    output [C_INPUT_FIFO_63_WIDTH-1:0] ap_fifo_iarg_63_dout,
    input ap_fifo_iarg_63_read,
    //input AXI-Stream to FIFO interface 64
    input s_axis_fifo_64_tlast,
    input s_axis_fifo_64_tvalid,
    input [C_INPUT_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tkeep,
    input [C_INPUT_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tstrb,
    input [C_INPUT_FIFO_64_DMWIDTH-1:0] s_axis_fifo_64_tdata,
    output s_axis_fifo_64_tready,
    output ap_fifo_iarg_64_empty_n,
    output [C_INPUT_FIFO_64_WIDTH-1:0] ap_fifo_iarg_64_dout,
    input ap_fifo_iarg_64_read,
    //input AXI-Stream to FIFO interface 65
    input s_axis_fifo_65_tlast,
    input s_axis_fifo_65_tvalid,
    input [C_INPUT_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tkeep,
    input [C_INPUT_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tstrb,
    input [C_INPUT_FIFO_65_DMWIDTH-1:0] s_axis_fifo_65_tdata,
    output s_axis_fifo_65_tready,
    output ap_fifo_iarg_65_empty_n,
    output [C_INPUT_FIFO_65_WIDTH-1:0] ap_fifo_iarg_65_dout,
    input ap_fifo_iarg_65_read,
    //input AXI-Stream to FIFO interface 66
    input s_axis_fifo_66_tlast,
    input s_axis_fifo_66_tvalid,
    input [C_INPUT_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tkeep,
    input [C_INPUT_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tstrb,
    input [C_INPUT_FIFO_66_DMWIDTH-1:0] s_axis_fifo_66_tdata,
    output s_axis_fifo_66_tready,
    output ap_fifo_iarg_66_empty_n,
    output [C_INPUT_FIFO_66_WIDTH-1:0] ap_fifo_iarg_66_dout,
    input ap_fifo_iarg_66_read,
    //input AXI-Stream to FIFO interface 67
    input s_axis_fifo_67_tlast,
    input s_axis_fifo_67_tvalid,
    input [C_INPUT_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tkeep,
    input [C_INPUT_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tstrb,
    input [C_INPUT_FIFO_67_DMWIDTH-1:0] s_axis_fifo_67_tdata,
    output s_axis_fifo_67_tready,
    output ap_fifo_iarg_67_empty_n,
    output [C_INPUT_FIFO_67_WIDTH-1:0] ap_fifo_iarg_67_dout,
    input ap_fifo_iarg_67_read,
    //input AXI-Stream to FIFO interface 68
    input s_axis_fifo_68_tlast,
    input s_axis_fifo_68_tvalid,
    input [C_INPUT_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tkeep,
    input [C_INPUT_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tstrb,
    input [C_INPUT_FIFO_68_DMWIDTH-1:0] s_axis_fifo_68_tdata,
    output s_axis_fifo_68_tready,
    output ap_fifo_iarg_68_empty_n,
    output [C_INPUT_FIFO_68_WIDTH-1:0] ap_fifo_iarg_68_dout,
    input ap_fifo_iarg_68_read,
    //input AXI-Stream to FIFO interface 69
    input s_axis_fifo_69_tlast,
    input s_axis_fifo_69_tvalid,
    input [C_INPUT_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tkeep,
    input [C_INPUT_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tstrb,
    input [C_INPUT_FIFO_69_DMWIDTH-1:0] s_axis_fifo_69_tdata,
    output s_axis_fifo_69_tready,
    output ap_fifo_iarg_69_empty_n,
    output [C_INPUT_FIFO_69_WIDTH-1:0] ap_fifo_iarg_69_dout,
    input ap_fifo_iarg_69_read,
    //input AXI-Stream to FIFO interface 70
    input s_axis_fifo_70_tlast,
    input s_axis_fifo_70_tvalid,
    input [C_INPUT_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tkeep,
    input [C_INPUT_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tstrb,
    input [C_INPUT_FIFO_70_DMWIDTH-1:0] s_axis_fifo_70_tdata,
    output s_axis_fifo_70_tready,
    output ap_fifo_iarg_70_empty_n,
    output [C_INPUT_FIFO_70_WIDTH-1:0] ap_fifo_iarg_70_dout,
    input ap_fifo_iarg_70_read,
    //input AXI-Stream to FIFO interface 71
    input s_axis_fifo_71_tlast,
    input s_axis_fifo_71_tvalid,
    input [C_INPUT_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tkeep,
    input [C_INPUT_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tstrb,
    input [C_INPUT_FIFO_71_DMWIDTH-1:0] s_axis_fifo_71_tdata,
    output s_axis_fifo_71_tready,
    output ap_fifo_iarg_71_empty_n,
    output [C_INPUT_FIFO_71_WIDTH-1:0] ap_fifo_iarg_71_dout,
    input ap_fifo_iarg_71_read,
    //input AXI-Stream to FIFO interface 72
    input s_axis_fifo_72_tlast,
    input s_axis_fifo_72_tvalid,
    input [C_INPUT_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tkeep,
    input [C_INPUT_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tstrb,
    input [C_INPUT_FIFO_72_DMWIDTH-1:0] s_axis_fifo_72_tdata,
    output s_axis_fifo_72_tready,
    output ap_fifo_iarg_72_empty_n,
    output [C_INPUT_FIFO_72_WIDTH-1:0] ap_fifo_iarg_72_dout,
    input ap_fifo_iarg_72_read,
    //input AXI-Stream to FIFO interface 73
    input s_axis_fifo_73_tlast,
    input s_axis_fifo_73_tvalid,
    input [C_INPUT_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tkeep,
    input [C_INPUT_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tstrb,
    input [C_INPUT_FIFO_73_DMWIDTH-1:0] s_axis_fifo_73_tdata,
    output s_axis_fifo_73_tready,
    output ap_fifo_iarg_73_empty_n,
    output [C_INPUT_FIFO_73_WIDTH-1:0] ap_fifo_iarg_73_dout,
    input ap_fifo_iarg_73_read,
    //input AXI-Stream to FIFO interface 74
    input s_axis_fifo_74_tlast,
    input s_axis_fifo_74_tvalid,
    input [C_INPUT_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tkeep,
    input [C_INPUT_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tstrb,
    input [C_INPUT_FIFO_74_DMWIDTH-1:0] s_axis_fifo_74_tdata,
    output s_axis_fifo_74_tready,
    output ap_fifo_iarg_74_empty_n,
    output [C_INPUT_FIFO_74_WIDTH-1:0] ap_fifo_iarg_74_dout,
    input ap_fifo_iarg_74_read,
    //input AXI-Stream to FIFO interface 75
    input s_axis_fifo_75_tlast,
    input s_axis_fifo_75_tvalid,
    input [C_INPUT_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tkeep,
    input [C_INPUT_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tstrb,
    input [C_INPUT_FIFO_75_DMWIDTH-1:0] s_axis_fifo_75_tdata,
    output s_axis_fifo_75_tready,
    output ap_fifo_iarg_75_empty_n,
    output [C_INPUT_FIFO_75_WIDTH-1:0] ap_fifo_iarg_75_dout,
    input ap_fifo_iarg_75_read,
    //input AXI-Stream to FIFO interface 76
    input s_axis_fifo_76_tlast,
    input s_axis_fifo_76_tvalid,
    input [C_INPUT_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tkeep,
    input [C_INPUT_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tstrb,
    input [C_INPUT_FIFO_76_DMWIDTH-1:0] s_axis_fifo_76_tdata,
    output s_axis_fifo_76_tready,
    output ap_fifo_iarg_76_empty_n,
    output [C_INPUT_FIFO_76_WIDTH-1:0] ap_fifo_iarg_76_dout,
    input ap_fifo_iarg_76_read,
    //input AXI-Stream to FIFO interface 77
    input s_axis_fifo_77_tlast,
    input s_axis_fifo_77_tvalid,
    input [C_INPUT_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tkeep,
    input [C_INPUT_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tstrb,
    input [C_INPUT_FIFO_77_DMWIDTH-1:0] s_axis_fifo_77_tdata,
    output s_axis_fifo_77_tready,
    output ap_fifo_iarg_77_empty_n,
    output [C_INPUT_FIFO_77_WIDTH-1:0] ap_fifo_iarg_77_dout,
    input ap_fifo_iarg_77_read,
    //input AXI-Stream to FIFO interface 78
    input s_axis_fifo_78_tlast,
    input s_axis_fifo_78_tvalid,
    input [C_INPUT_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tkeep,
    input [C_INPUT_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tstrb,
    input [C_INPUT_FIFO_78_DMWIDTH-1:0] s_axis_fifo_78_tdata,
    output s_axis_fifo_78_tready,
    output ap_fifo_iarg_78_empty_n,
    output [C_INPUT_FIFO_78_WIDTH-1:0] ap_fifo_iarg_78_dout,
    input ap_fifo_iarg_78_read,
    //input AXI-Stream to FIFO interface 79
    input s_axis_fifo_79_tlast,
    input s_axis_fifo_79_tvalid,
    input [C_INPUT_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tkeep,
    input [C_INPUT_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tstrb,
    input [C_INPUT_FIFO_79_DMWIDTH-1:0] s_axis_fifo_79_tdata,
    output s_axis_fifo_79_tready,
    output ap_fifo_iarg_79_empty_n,
    output [C_INPUT_FIFO_79_WIDTH-1:0] ap_fifo_iarg_79_dout,
    input ap_fifo_iarg_79_read,
    //input AXI-Stream to FIFO interface 80
    input s_axis_fifo_80_tlast,
    input s_axis_fifo_80_tvalid,
    input [C_INPUT_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tkeep,
    input [C_INPUT_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tstrb,
    input [C_INPUT_FIFO_80_DMWIDTH-1:0] s_axis_fifo_80_tdata,
    output s_axis_fifo_80_tready,
    output ap_fifo_iarg_80_empty_n,
    output [C_INPUT_FIFO_80_WIDTH-1:0] ap_fifo_iarg_80_dout,
    input ap_fifo_iarg_80_read,
    //input AXI-Stream to FIFO interface 81
    input s_axis_fifo_81_tlast,
    input s_axis_fifo_81_tvalid,
    input [C_INPUT_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tkeep,
    input [C_INPUT_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tstrb,
    input [C_INPUT_FIFO_81_DMWIDTH-1:0] s_axis_fifo_81_tdata,
    output s_axis_fifo_81_tready,
    output ap_fifo_iarg_81_empty_n,
    output [C_INPUT_FIFO_81_WIDTH-1:0] ap_fifo_iarg_81_dout,
    input ap_fifo_iarg_81_read,
    //input AXI-Stream to FIFO interface 82
    input s_axis_fifo_82_tlast,
    input s_axis_fifo_82_tvalid,
    input [C_INPUT_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tkeep,
    input [C_INPUT_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tstrb,
    input [C_INPUT_FIFO_82_DMWIDTH-1:0] s_axis_fifo_82_tdata,
    output s_axis_fifo_82_tready,
    output ap_fifo_iarg_82_empty_n,
    output [C_INPUT_FIFO_82_WIDTH-1:0] ap_fifo_iarg_82_dout,
    input ap_fifo_iarg_82_read,
    //input AXI-Stream to FIFO interface 83
    input s_axis_fifo_83_tlast,
    input s_axis_fifo_83_tvalid,
    input [C_INPUT_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tkeep,
    input [C_INPUT_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tstrb,
    input [C_INPUT_FIFO_83_DMWIDTH-1:0] s_axis_fifo_83_tdata,
    output s_axis_fifo_83_tready,
    output ap_fifo_iarg_83_empty_n,
    output [C_INPUT_FIFO_83_WIDTH-1:0] ap_fifo_iarg_83_dout,
    input ap_fifo_iarg_83_read,
    //input AXI-Stream to FIFO interface 84
    input s_axis_fifo_84_tlast,
    input s_axis_fifo_84_tvalid,
    input [C_INPUT_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tkeep,
    input [C_INPUT_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tstrb,
    input [C_INPUT_FIFO_84_DMWIDTH-1:0] s_axis_fifo_84_tdata,
    output s_axis_fifo_84_tready,
    output ap_fifo_iarg_84_empty_n,
    output [C_INPUT_FIFO_84_WIDTH-1:0] ap_fifo_iarg_84_dout,
    input ap_fifo_iarg_84_read,
    //input AXI-Stream to FIFO interface 85
    input s_axis_fifo_85_tlast,
    input s_axis_fifo_85_tvalid,
    input [C_INPUT_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tkeep,
    input [C_INPUT_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tstrb,
    input [C_INPUT_FIFO_85_DMWIDTH-1:0] s_axis_fifo_85_tdata,
    output s_axis_fifo_85_tready,
    output ap_fifo_iarg_85_empty_n,
    output [C_INPUT_FIFO_85_WIDTH-1:0] ap_fifo_iarg_85_dout,
    input ap_fifo_iarg_85_read,
    //input AXI-Stream to FIFO interface 86
    input s_axis_fifo_86_tlast,
    input s_axis_fifo_86_tvalid,
    input [C_INPUT_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tkeep,
    input [C_INPUT_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tstrb,
    input [C_INPUT_FIFO_86_DMWIDTH-1:0] s_axis_fifo_86_tdata,
    output s_axis_fifo_86_tready,
    output ap_fifo_iarg_86_empty_n,
    output [C_INPUT_FIFO_86_WIDTH-1:0] ap_fifo_iarg_86_dout,
    input ap_fifo_iarg_86_read,
    //input AXI-Stream to FIFO interface 87
    input s_axis_fifo_87_tlast,
    input s_axis_fifo_87_tvalid,
    input [C_INPUT_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tkeep,
    input [C_INPUT_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tstrb,
    input [C_INPUT_FIFO_87_DMWIDTH-1:0] s_axis_fifo_87_tdata,
    output s_axis_fifo_87_tready,
    output ap_fifo_iarg_87_empty_n,
    output [C_INPUT_FIFO_87_WIDTH-1:0] ap_fifo_iarg_87_dout,
    input ap_fifo_iarg_87_read,
    //input AXI-Stream to FIFO interface 88
    input s_axis_fifo_88_tlast,
    input s_axis_fifo_88_tvalid,
    input [C_INPUT_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tkeep,
    input [C_INPUT_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tstrb,
    input [C_INPUT_FIFO_88_DMWIDTH-1:0] s_axis_fifo_88_tdata,
    output s_axis_fifo_88_tready,
    output ap_fifo_iarg_88_empty_n,
    output [C_INPUT_FIFO_88_WIDTH-1:0] ap_fifo_iarg_88_dout,
    input ap_fifo_iarg_88_read,
    //input AXI-Stream to FIFO interface 89
    input s_axis_fifo_89_tlast,
    input s_axis_fifo_89_tvalid,
    input [C_INPUT_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tkeep,
    input [C_INPUT_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tstrb,
    input [C_INPUT_FIFO_89_DMWIDTH-1:0] s_axis_fifo_89_tdata,
    output s_axis_fifo_89_tready,
    output ap_fifo_iarg_89_empty_n,
    output [C_INPUT_FIFO_89_WIDTH-1:0] ap_fifo_iarg_89_dout,
    input ap_fifo_iarg_89_read,
    //input AXI-Stream to FIFO interface 90
    input s_axis_fifo_90_tlast,
    input s_axis_fifo_90_tvalid,
    input [C_INPUT_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tkeep,
    input [C_INPUT_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tstrb,
    input [C_INPUT_FIFO_90_DMWIDTH-1:0] s_axis_fifo_90_tdata,
    output s_axis_fifo_90_tready,
    output ap_fifo_iarg_90_empty_n,
    output [C_INPUT_FIFO_90_WIDTH-1:0] ap_fifo_iarg_90_dout,
    input ap_fifo_iarg_90_read,
    //input AXI-Stream to FIFO interface 91
    input s_axis_fifo_91_tlast,
    input s_axis_fifo_91_tvalid,
    input [C_INPUT_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tkeep,
    input [C_INPUT_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tstrb,
    input [C_INPUT_FIFO_91_DMWIDTH-1:0] s_axis_fifo_91_tdata,
    output s_axis_fifo_91_tready,
    output ap_fifo_iarg_91_empty_n,
    output [C_INPUT_FIFO_91_WIDTH-1:0] ap_fifo_iarg_91_dout,
    input ap_fifo_iarg_91_read,
    //input AXI-Stream to FIFO interface 92
    input s_axis_fifo_92_tlast,
    input s_axis_fifo_92_tvalid,
    input [C_INPUT_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tkeep,
    input [C_INPUT_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tstrb,
    input [C_INPUT_FIFO_92_DMWIDTH-1:0] s_axis_fifo_92_tdata,
    output s_axis_fifo_92_tready,
    output ap_fifo_iarg_92_empty_n,
    output [C_INPUT_FIFO_92_WIDTH-1:0] ap_fifo_iarg_92_dout,
    input ap_fifo_iarg_92_read,
    //input AXI-Stream to FIFO interface 93
    input s_axis_fifo_93_tlast,
    input s_axis_fifo_93_tvalid,
    input [C_INPUT_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tkeep,
    input [C_INPUT_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tstrb,
    input [C_INPUT_FIFO_93_DMWIDTH-1:0] s_axis_fifo_93_tdata,
    output s_axis_fifo_93_tready,
    output ap_fifo_iarg_93_empty_n,
    output [C_INPUT_FIFO_93_WIDTH-1:0] ap_fifo_iarg_93_dout,
    input ap_fifo_iarg_93_read,
    //input AXI-Stream to FIFO interface 94
    input s_axis_fifo_94_tlast,
    input s_axis_fifo_94_tvalid,
    input [C_INPUT_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tkeep,
    input [C_INPUT_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tstrb,
    input [C_INPUT_FIFO_94_DMWIDTH-1:0] s_axis_fifo_94_tdata,
    output s_axis_fifo_94_tready,
    output ap_fifo_iarg_94_empty_n,
    output [C_INPUT_FIFO_94_WIDTH-1:0] ap_fifo_iarg_94_dout,
    input ap_fifo_iarg_94_read,
    //input AXI-Stream to FIFO interface 95
    input s_axis_fifo_95_tlast,
    input s_axis_fifo_95_tvalid,
    input [C_INPUT_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tkeep,
    input [C_INPUT_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tstrb,
    input [C_INPUT_FIFO_95_DMWIDTH-1:0] s_axis_fifo_95_tdata,
    output s_axis_fifo_95_tready,
    output ap_fifo_iarg_95_empty_n,
    output [C_INPUT_FIFO_95_WIDTH-1:0] ap_fifo_iarg_95_dout,
    input ap_fifo_iarg_95_read,
    //input AXI-Stream to FIFO interface 96
    input s_axis_fifo_96_tlast,
    input s_axis_fifo_96_tvalid,
    input [C_INPUT_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tkeep,
    input [C_INPUT_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tstrb,
    input [C_INPUT_FIFO_96_DMWIDTH-1:0] s_axis_fifo_96_tdata,
    output s_axis_fifo_96_tready,
    output ap_fifo_iarg_96_empty_n,
    output [C_INPUT_FIFO_96_WIDTH-1:0] ap_fifo_iarg_96_dout,
    input ap_fifo_iarg_96_read,
    //input AXI-Stream to FIFO interface 97
    input s_axis_fifo_97_tlast,
    input s_axis_fifo_97_tvalid,
    input [C_INPUT_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tkeep,
    input [C_INPUT_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tstrb,
    input [C_INPUT_FIFO_97_DMWIDTH-1:0] s_axis_fifo_97_tdata,
    output s_axis_fifo_97_tready,
    output ap_fifo_iarg_97_empty_n,
    output [C_INPUT_FIFO_97_WIDTH-1:0] ap_fifo_iarg_97_dout,
    input ap_fifo_iarg_97_read,
    //input AXI-Stream to FIFO interface 98
    input s_axis_fifo_98_tlast,
    input s_axis_fifo_98_tvalid,
    input [C_INPUT_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tkeep,
    input [C_INPUT_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tstrb,
    input [C_INPUT_FIFO_98_DMWIDTH-1:0] s_axis_fifo_98_tdata,
    output s_axis_fifo_98_tready,
    output ap_fifo_iarg_98_empty_n,
    output [C_INPUT_FIFO_98_WIDTH-1:0] ap_fifo_iarg_98_dout,
    input ap_fifo_iarg_98_read,
    //input AXI-Stream to FIFO interface 99
    input s_axis_fifo_99_tlast,
    input s_axis_fifo_99_tvalid,
    input [C_INPUT_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tkeep,
    input [C_INPUT_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tstrb,
    input [C_INPUT_FIFO_99_DMWIDTH-1:0] s_axis_fifo_99_tdata,
    output s_axis_fifo_99_tready,
    output ap_fifo_iarg_99_empty_n,
    output [C_INPUT_FIFO_99_WIDTH-1:0] ap_fifo_iarg_99_dout,
    input ap_fifo_iarg_99_read,
    //input AXI-Stream to FIFO interface 100
    input s_axis_fifo_100_tlast,
    input s_axis_fifo_100_tvalid,
    input [C_INPUT_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tkeep,
    input [C_INPUT_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tstrb,
    input [C_INPUT_FIFO_100_DMWIDTH-1:0] s_axis_fifo_100_tdata,
    output s_axis_fifo_100_tready,
    output ap_fifo_iarg_100_empty_n,
    output [C_INPUT_FIFO_100_WIDTH-1:0] ap_fifo_iarg_100_dout,
    input ap_fifo_iarg_100_read,
    //input AXI-Stream to FIFO interface 101
    input s_axis_fifo_101_tlast,
    input s_axis_fifo_101_tvalid,
    input [C_INPUT_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tkeep,
    input [C_INPUT_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tstrb,
    input [C_INPUT_FIFO_101_DMWIDTH-1:0] s_axis_fifo_101_tdata,
    output s_axis_fifo_101_tready,
    output ap_fifo_iarg_101_empty_n,
    output [C_INPUT_FIFO_101_WIDTH-1:0] ap_fifo_iarg_101_dout,
    input ap_fifo_iarg_101_read,
    //input AXI-Stream to FIFO interface 102
    input s_axis_fifo_102_tlast,
    input s_axis_fifo_102_tvalid,
    input [C_INPUT_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tkeep,
    input [C_INPUT_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tstrb,
    input [C_INPUT_FIFO_102_DMWIDTH-1:0] s_axis_fifo_102_tdata,
    output s_axis_fifo_102_tready,
    output ap_fifo_iarg_102_empty_n,
    output [C_INPUT_FIFO_102_WIDTH-1:0] ap_fifo_iarg_102_dout,
    input ap_fifo_iarg_102_read,
    //input AXI-Stream to FIFO interface 103
    input s_axis_fifo_103_tlast,
    input s_axis_fifo_103_tvalid,
    input [C_INPUT_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tkeep,
    input [C_INPUT_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tstrb,
    input [C_INPUT_FIFO_103_DMWIDTH-1:0] s_axis_fifo_103_tdata,
    output s_axis_fifo_103_tready,
    output ap_fifo_iarg_103_empty_n,
    output [C_INPUT_FIFO_103_WIDTH-1:0] ap_fifo_iarg_103_dout,
    input ap_fifo_iarg_103_read,
    //input AXI-Stream to FIFO interface 104
    input s_axis_fifo_104_tlast,
    input s_axis_fifo_104_tvalid,
    input [C_INPUT_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tkeep,
    input [C_INPUT_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tstrb,
    input [C_INPUT_FIFO_104_DMWIDTH-1:0] s_axis_fifo_104_tdata,
    output s_axis_fifo_104_tready,
    output ap_fifo_iarg_104_empty_n,
    output [C_INPUT_FIFO_104_WIDTH-1:0] ap_fifo_iarg_104_dout,
    input ap_fifo_iarg_104_read,
    //input AXI-Stream to FIFO interface 105
    input s_axis_fifo_105_tlast,
    input s_axis_fifo_105_tvalid,
    input [C_INPUT_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tkeep,
    input [C_INPUT_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tstrb,
    input [C_INPUT_FIFO_105_DMWIDTH-1:0] s_axis_fifo_105_tdata,
    output s_axis_fifo_105_tready,
    output ap_fifo_iarg_105_empty_n,
    output [C_INPUT_FIFO_105_WIDTH-1:0] ap_fifo_iarg_105_dout,
    input ap_fifo_iarg_105_read,
    //input AXI-Stream to FIFO interface 106
    input s_axis_fifo_106_tlast,
    input s_axis_fifo_106_tvalid,
    input [C_INPUT_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tkeep,
    input [C_INPUT_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tstrb,
    input [C_INPUT_FIFO_106_DMWIDTH-1:0] s_axis_fifo_106_tdata,
    output s_axis_fifo_106_tready,
    output ap_fifo_iarg_106_empty_n,
    output [C_INPUT_FIFO_106_WIDTH-1:0] ap_fifo_iarg_106_dout,
    input ap_fifo_iarg_106_read,
    //input AXI-Stream to FIFO interface 107
    input s_axis_fifo_107_tlast,
    input s_axis_fifo_107_tvalid,
    input [C_INPUT_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tkeep,
    input [C_INPUT_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tstrb,
    input [C_INPUT_FIFO_107_DMWIDTH-1:0] s_axis_fifo_107_tdata,
    output s_axis_fifo_107_tready,
    output ap_fifo_iarg_107_empty_n,
    output [C_INPUT_FIFO_107_WIDTH-1:0] ap_fifo_iarg_107_dout,
    input ap_fifo_iarg_107_read,
    //input AXI-Stream to FIFO interface 108
    input s_axis_fifo_108_tlast,
    input s_axis_fifo_108_tvalid,
    input [C_INPUT_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tkeep,
    input [C_INPUT_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tstrb,
    input [C_INPUT_FIFO_108_DMWIDTH-1:0] s_axis_fifo_108_tdata,
    output s_axis_fifo_108_tready,
    output ap_fifo_iarg_108_empty_n,
    output [C_INPUT_FIFO_108_WIDTH-1:0] ap_fifo_iarg_108_dout,
    input ap_fifo_iarg_108_read,
    //input AXI-Stream to FIFO interface 109
    input s_axis_fifo_109_tlast,
    input s_axis_fifo_109_tvalid,
    input [C_INPUT_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tkeep,
    input [C_INPUT_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tstrb,
    input [C_INPUT_FIFO_109_DMWIDTH-1:0] s_axis_fifo_109_tdata,
    output s_axis_fifo_109_tready,
    output ap_fifo_iarg_109_empty_n,
    output [C_INPUT_FIFO_109_WIDTH-1:0] ap_fifo_iarg_109_dout,
    input ap_fifo_iarg_109_read,
    //input AXI-Stream to FIFO interface 110
    input s_axis_fifo_110_tlast,
    input s_axis_fifo_110_tvalid,
    input [C_INPUT_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tkeep,
    input [C_INPUT_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tstrb,
    input [C_INPUT_FIFO_110_DMWIDTH-1:0] s_axis_fifo_110_tdata,
    output s_axis_fifo_110_tready,
    output ap_fifo_iarg_110_empty_n,
    output [C_INPUT_FIFO_110_WIDTH-1:0] ap_fifo_iarg_110_dout,
    input ap_fifo_iarg_110_read,
    //input AXI-Stream to FIFO interface 111
    input s_axis_fifo_111_tlast,
    input s_axis_fifo_111_tvalid,
    input [C_INPUT_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tkeep,
    input [C_INPUT_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tstrb,
    input [C_INPUT_FIFO_111_DMWIDTH-1:0] s_axis_fifo_111_tdata,
    output s_axis_fifo_111_tready,
    output ap_fifo_iarg_111_empty_n,
    output [C_INPUT_FIFO_111_WIDTH-1:0] ap_fifo_iarg_111_dout,
    input ap_fifo_iarg_111_read,
    //input AXI-Stream to FIFO interface 112
    input s_axis_fifo_112_tlast,
    input s_axis_fifo_112_tvalid,
    input [C_INPUT_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tkeep,
    input [C_INPUT_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tstrb,
    input [C_INPUT_FIFO_112_DMWIDTH-1:0] s_axis_fifo_112_tdata,
    output s_axis_fifo_112_tready,
    output ap_fifo_iarg_112_empty_n,
    output [C_INPUT_FIFO_112_WIDTH-1:0] ap_fifo_iarg_112_dout,
    input ap_fifo_iarg_112_read,
    //input AXI-Stream to FIFO interface 113
    input s_axis_fifo_113_tlast,
    input s_axis_fifo_113_tvalid,
    input [C_INPUT_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tkeep,
    input [C_INPUT_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tstrb,
    input [C_INPUT_FIFO_113_DMWIDTH-1:0] s_axis_fifo_113_tdata,
    output s_axis_fifo_113_tready,
    output ap_fifo_iarg_113_empty_n,
    output [C_INPUT_FIFO_113_WIDTH-1:0] ap_fifo_iarg_113_dout,
    input ap_fifo_iarg_113_read,
    //input AXI-Stream to FIFO interface 114
    input s_axis_fifo_114_tlast,
    input s_axis_fifo_114_tvalid,
    input [C_INPUT_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tkeep,
    input [C_INPUT_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tstrb,
    input [C_INPUT_FIFO_114_DMWIDTH-1:0] s_axis_fifo_114_tdata,
    output s_axis_fifo_114_tready,
    output ap_fifo_iarg_114_empty_n,
    output [C_INPUT_FIFO_114_WIDTH-1:0] ap_fifo_iarg_114_dout,
    input ap_fifo_iarg_114_read,
    //input AXI-Stream to FIFO interface 115
    input s_axis_fifo_115_tlast,
    input s_axis_fifo_115_tvalid,
    input [C_INPUT_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tkeep,
    input [C_INPUT_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tstrb,
    input [C_INPUT_FIFO_115_DMWIDTH-1:0] s_axis_fifo_115_tdata,
    output s_axis_fifo_115_tready,
    output ap_fifo_iarg_115_empty_n,
    output [C_INPUT_FIFO_115_WIDTH-1:0] ap_fifo_iarg_115_dout,
    input ap_fifo_iarg_115_read,
    //input AXI-Stream to FIFO interface 116
    input s_axis_fifo_116_tlast,
    input s_axis_fifo_116_tvalid,
    input [C_INPUT_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tkeep,
    input [C_INPUT_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tstrb,
    input [C_INPUT_FIFO_116_DMWIDTH-1:0] s_axis_fifo_116_tdata,
    output s_axis_fifo_116_tready,
    output ap_fifo_iarg_116_empty_n,
    output [C_INPUT_FIFO_116_WIDTH-1:0] ap_fifo_iarg_116_dout,
    input ap_fifo_iarg_116_read,
    //input AXI-Stream to FIFO interface 117
    input s_axis_fifo_117_tlast,
    input s_axis_fifo_117_tvalid,
    input [C_INPUT_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tkeep,
    input [C_INPUT_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tstrb,
    input [C_INPUT_FIFO_117_DMWIDTH-1:0] s_axis_fifo_117_tdata,
    output s_axis_fifo_117_tready,
    output ap_fifo_iarg_117_empty_n,
    output [C_INPUT_FIFO_117_WIDTH-1:0] ap_fifo_iarg_117_dout,
    input ap_fifo_iarg_117_read,
    //input AXI-Stream to FIFO interface 118
    input s_axis_fifo_118_tlast,
    input s_axis_fifo_118_tvalid,
    input [C_INPUT_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tkeep,
    input [C_INPUT_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tstrb,
    input [C_INPUT_FIFO_118_DMWIDTH-1:0] s_axis_fifo_118_tdata,
    output s_axis_fifo_118_tready,
    output ap_fifo_iarg_118_empty_n,
    output [C_INPUT_FIFO_118_WIDTH-1:0] ap_fifo_iarg_118_dout,
    input ap_fifo_iarg_118_read,
    //input AXI-Stream to FIFO interface 119
    input s_axis_fifo_119_tlast,
    input s_axis_fifo_119_tvalid,
    input [C_INPUT_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tkeep,
    input [C_INPUT_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tstrb,
    input [C_INPUT_FIFO_119_DMWIDTH-1:0] s_axis_fifo_119_tdata,
    output s_axis_fifo_119_tready,
    output ap_fifo_iarg_119_empty_n,
    output [C_INPUT_FIFO_119_WIDTH-1:0] ap_fifo_iarg_119_dout,
    input ap_fifo_iarg_119_read,
    //input AXI-Stream to FIFO interface 120
    input s_axis_fifo_120_tlast,
    input s_axis_fifo_120_tvalid,
    input [C_INPUT_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tkeep,
    input [C_INPUT_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tstrb,
    input [C_INPUT_FIFO_120_DMWIDTH-1:0] s_axis_fifo_120_tdata,
    output s_axis_fifo_120_tready,
    output ap_fifo_iarg_120_empty_n,
    output [C_INPUT_FIFO_120_WIDTH-1:0] ap_fifo_iarg_120_dout,
    input ap_fifo_iarg_120_read,
    //input AXI-Stream to FIFO interface 121
    input s_axis_fifo_121_tlast,
    input s_axis_fifo_121_tvalid,
    input [C_INPUT_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tkeep,
    input [C_INPUT_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tstrb,
    input [C_INPUT_FIFO_121_DMWIDTH-1:0] s_axis_fifo_121_tdata,
    output s_axis_fifo_121_tready,
    output ap_fifo_iarg_121_empty_n,
    output [C_INPUT_FIFO_121_WIDTH-1:0] ap_fifo_iarg_121_dout,
    input ap_fifo_iarg_121_read,
    //input AXI-Stream to FIFO interface 122
    input s_axis_fifo_122_tlast,
    input s_axis_fifo_122_tvalid,
    input [C_INPUT_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tkeep,
    input [C_INPUT_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tstrb,
    input [C_INPUT_FIFO_122_DMWIDTH-1:0] s_axis_fifo_122_tdata,
    output s_axis_fifo_122_tready,
    output ap_fifo_iarg_122_empty_n,
    output [C_INPUT_FIFO_122_WIDTH-1:0] ap_fifo_iarg_122_dout,
    input ap_fifo_iarg_122_read,
    //input AXI-Stream to FIFO interface 123
    input s_axis_fifo_123_tlast,
    input s_axis_fifo_123_tvalid,
    input [C_INPUT_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tkeep,
    input [C_INPUT_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tstrb,
    input [C_INPUT_FIFO_123_DMWIDTH-1:0] s_axis_fifo_123_tdata,
    output s_axis_fifo_123_tready,
    output ap_fifo_iarg_123_empty_n,
    output [C_INPUT_FIFO_123_WIDTH-1:0] ap_fifo_iarg_123_dout,
    input ap_fifo_iarg_123_read,
    //input AXI-Stream to FIFO interface 124
    input s_axis_fifo_124_tlast,
    input s_axis_fifo_124_tvalid,
    input [C_INPUT_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tkeep,
    input [C_INPUT_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tstrb,
    input [C_INPUT_FIFO_124_DMWIDTH-1:0] s_axis_fifo_124_tdata,
    output s_axis_fifo_124_tready,
    output ap_fifo_iarg_124_empty_n,
    output [C_INPUT_FIFO_124_WIDTH-1:0] ap_fifo_iarg_124_dout,
    input ap_fifo_iarg_124_read,
    //input AXI-Stream to FIFO interface 125
    input s_axis_fifo_125_tlast,
    input s_axis_fifo_125_tvalid,
    input [C_INPUT_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tkeep,
    input [C_INPUT_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tstrb,
    input [C_INPUT_FIFO_125_DMWIDTH-1:0] s_axis_fifo_125_tdata,
    output s_axis_fifo_125_tready,
    output ap_fifo_iarg_125_empty_n,
    output [C_INPUT_FIFO_125_WIDTH-1:0] ap_fifo_iarg_125_dout,
    input ap_fifo_iarg_125_read,
    //input AXI-Stream to FIFO interface 126
    input s_axis_fifo_126_tlast,
    input s_axis_fifo_126_tvalid,
    input [C_INPUT_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tkeep,
    input [C_INPUT_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tstrb,
    input [C_INPUT_FIFO_126_DMWIDTH-1:0] s_axis_fifo_126_tdata,
    output s_axis_fifo_126_tready,
    output ap_fifo_iarg_126_empty_n,
    output [C_INPUT_FIFO_126_WIDTH-1:0] ap_fifo_iarg_126_dout,
    input ap_fifo_iarg_126_read,
    //input AXI-Stream to FIFO interface 127
    input s_axis_fifo_127_tlast,
    input s_axis_fifo_127_tvalid,
    input [C_INPUT_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tkeep,
    input [C_INPUT_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tstrb,
    input [C_INPUT_FIFO_127_DMWIDTH-1:0] s_axis_fifo_127_tdata,
    output s_axis_fifo_127_tready,
    output ap_fifo_iarg_127_empty_n,
    output [C_INPUT_FIFO_127_WIDTH-1:0] ap_fifo_iarg_127_dout,
    input ap_fifo_iarg_127_read,
    //-----------------------------------------------------
    //output FIFO to AXI-Stream interface 0
    output m_axis_fifo_0_tlast,
    output m_axis_fifo_0_tvalid,
    output [C_OUTPUT_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tkeep,
    output [C_OUTPUT_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tstrb,
    output [C_OUTPUT_FIFO_0_DMWIDTH-1:0] m_axis_fifo_0_tdata,
    input m_axis_fifo_0_tready,
    output ap_fifo_oarg_0_full_n,
    input [C_OUTPUT_FIFO_0_WIDTH-1:0] ap_fifo_oarg_0_din,
    input ap_fifo_oarg_0_write,
    //output FIFO to AXI-Stream interface 1
    output m_axis_fifo_1_tlast,
    output m_axis_fifo_1_tvalid,
    output [C_OUTPUT_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tkeep,
    output [C_OUTPUT_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tstrb,
    output [C_OUTPUT_FIFO_1_DMWIDTH-1:0] m_axis_fifo_1_tdata,
    input m_axis_fifo_1_tready,
    output ap_fifo_oarg_1_full_n,
    input [C_OUTPUT_FIFO_1_WIDTH-1:0] ap_fifo_oarg_1_din,
    input ap_fifo_oarg_1_write,
    //output FIFO to AXI-Stream interface 2
    output m_axis_fifo_2_tlast,
    output m_axis_fifo_2_tvalid,
    output [C_OUTPUT_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tkeep,
    output [C_OUTPUT_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tstrb,
    output [C_OUTPUT_FIFO_2_DMWIDTH-1:0] m_axis_fifo_2_tdata,
    input m_axis_fifo_2_tready,
    output ap_fifo_oarg_2_full_n,
    input [C_OUTPUT_FIFO_2_WIDTH-1:0] ap_fifo_oarg_2_din,
    input ap_fifo_oarg_2_write,
    //output FIFO to AXI-Stream interface 3
    output m_axis_fifo_3_tlast,
    output m_axis_fifo_3_tvalid,
    output [C_OUTPUT_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tkeep,
    output [C_OUTPUT_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tstrb,
    output [C_OUTPUT_FIFO_3_DMWIDTH-1:0] m_axis_fifo_3_tdata,
    input m_axis_fifo_3_tready,
    output ap_fifo_oarg_3_full_n,
    input [C_OUTPUT_FIFO_3_WIDTH-1:0] ap_fifo_oarg_3_din,
    input ap_fifo_oarg_3_write,
    //output FIFO to AXI-Stream interface 4
    output m_axis_fifo_4_tlast,
    output m_axis_fifo_4_tvalid,
    output [C_OUTPUT_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tkeep,
    output [C_OUTPUT_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tstrb,
    output [C_OUTPUT_FIFO_4_DMWIDTH-1:0] m_axis_fifo_4_tdata,
    input m_axis_fifo_4_tready,
    output ap_fifo_oarg_4_full_n,
    input [C_OUTPUT_FIFO_4_WIDTH-1:0] ap_fifo_oarg_4_din,
    input ap_fifo_oarg_4_write,
    //output FIFO to AXI-Stream interface 5
    output m_axis_fifo_5_tlast,
    output m_axis_fifo_5_tvalid,
    output [C_OUTPUT_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tkeep,
    output [C_OUTPUT_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tstrb,
    output [C_OUTPUT_FIFO_5_DMWIDTH-1:0] m_axis_fifo_5_tdata,
    input m_axis_fifo_5_tready,
    output ap_fifo_oarg_5_full_n,
    input [C_OUTPUT_FIFO_5_WIDTH-1:0] ap_fifo_oarg_5_din,
    input ap_fifo_oarg_5_write,
    //output FIFO to AXI-Stream interface 6
    output m_axis_fifo_6_tlast,
    output m_axis_fifo_6_tvalid,
    output [C_OUTPUT_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tkeep,
    output [C_OUTPUT_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tstrb,
    output [C_OUTPUT_FIFO_6_DMWIDTH-1:0] m_axis_fifo_6_tdata,
    input m_axis_fifo_6_tready,
    output ap_fifo_oarg_6_full_n,
    input [C_OUTPUT_FIFO_6_WIDTH-1:0] ap_fifo_oarg_6_din,
    input ap_fifo_oarg_6_write,
    //output FIFO to AXI-Stream interface 7
    output m_axis_fifo_7_tlast,
    output m_axis_fifo_7_tvalid,
    output [C_OUTPUT_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tkeep,
    output [C_OUTPUT_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tstrb,
    output [C_OUTPUT_FIFO_7_DMWIDTH-1:0] m_axis_fifo_7_tdata,
    input m_axis_fifo_7_tready,
    output ap_fifo_oarg_7_full_n,
    input [C_OUTPUT_FIFO_7_WIDTH-1:0] ap_fifo_oarg_7_din,
    input ap_fifo_oarg_7_write,
    //output FIFO to AXI-Stream interface 8
    output m_axis_fifo_8_tlast,
    output m_axis_fifo_8_tvalid,
    output [C_OUTPUT_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tkeep,
    output [C_OUTPUT_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tstrb,
    output [C_OUTPUT_FIFO_8_DMWIDTH-1:0] m_axis_fifo_8_tdata,
    input m_axis_fifo_8_tready,
    output ap_fifo_oarg_8_full_n,
    input [C_OUTPUT_FIFO_8_WIDTH-1:0] ap_fifo_oarg_8_din,
    input ap_fifo_oarg_8_write,
    //output FIFO to AXI-Stream interface 9
    output m_axis_fifo_9_tlast,
    output m_axis_fifo_9_tvalid,
    output [C_OUTPUT_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tkeep,
    output [C_OUTPUT_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tstrb,
    output [C_OUTPUT_FIFO_9_DMWIDTH-1:0] m_axis_fifo_9_tdata,
    input m_axis_fifo_9_tready,
    output ap_fifo_oarg_9_full_n,
    input [C_OUTPUT_FIFO_9_WIDTH-1:0] ap_fifo_oarg_9_din,
    input ap_fifo_oarg_9_write,
    //output FIFO to AXI-Stream interface 10
    output m_axis_fifo_10_tlast,
    output m_axis_fifo_10_tvalid,
    output [C_OUTPUT_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tkeep,
    output [C_OUTPUT_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tstrb,
    output [C_OUTPUT_FIFO_10_DMWIDTH-1:0] m_axis_fifo_10_tdata,
    input m_axis_fifo_10_tready,
    output ap_fifo_oarg_10_full_n,
    input [C_OUTPUT_FIFO_10_WIDTH-1:0] ap_fifo_oarg_10_din,
    input ap_fifo_oarg_10_write,
    //output FIFO to AXI-Stream interface 11
    output m_axis_fifo_11_tlast,
    output m_axis_fifo_11_tvalid,
    output [C_OUTPUT_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tkeep,
    output [C_OUTPUT_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tstrb,
    output [C_OUTPUT_FIFO_11_DMWIDTH-1:0] m_axis_fifo_11_tdata,
    input m_axis_fifo_11_tready,
    output ap_fifo_oarg_11_full_n,
    input [C_OUTPUT_FIFO_11_WIDTH-1:0] ap_fifo_oarg_11_din,
    input ap_fifo_oarg_11_write,
    //output FIFO to AXI-Stream interface 12
    output m_axis_fifo_12_tlast,
    output m_axis_fifo_12_tvalid,
    output [C_OUTPUT_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tkeep,
    output [C_OUTPUT_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tstrb,
    output [C_OUTPUT_FIFO_12_DMWIDTH-1:0] m_axis_fifo_12_tdata,
    input m_axis_fifo_12_tready,
    output ap_fifo_oarg_12_full_n,
    input [C_OUTPUT_FIFO_12_WIDTH-1:0] ap_fifo_oarg_12_din,
    input ap_fifo_oarg_12_write,
    //output FIFO to AXI-Stream interface 13
    output m_axis_fifo_13_tlast,
    output m_axis_fifo_13_tvalid,
    output [C_OUTPUT_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tkeep,
    output [C_OUTPUT_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tstrb,
    output [C_OUTPUT_FIFO_13_DMWIDTH-1:0] m_axis_fifo_13_tdata,
    input m_axis_fifo_13_tready,
    output ap_fifo_oarg_13_full_n,
    input [C_OUTPUT_FIFO_13_WIDTH-1:0] ap_fifo_oarg_13_din,
    input ap_fifo_oarg_13_write,
    //output FIFO to AXI-Stream interface 14
    output m_axis_fifo_14_tlast,
    output m_axis_fifo_14_tvalid,
    output [C_OUTPUT_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tkeep,
    output [C_OUTPUT_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tstrb,
    output [C_OUTPUT_FIFO_14_DMWIDTH-1:0] m_axis_fifo_14_tdata,
    input m_axis_fifo_14_tready,
    output ap_fifo_oarg_14_full_n,
    input [C_OUTPUT_FIFO_14_WIDTH-1:0] ap_fifo_oarg_14_din,
    input ap_fifo_oarg_14_write,
    //output FIFO to AXI-Stream interface 15
    output m_axis_fifo_15_tlast,
    output m_axis_fifo_15_tvalid,
    output [C_OUTPUT_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tkeep,
    output [C_OUTPUT_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tstrb,
    output [C_OUTPUT_FIFO_15_DMWIDTH-1:0] m_axis_fifo_15_tdata,
    input m_axis_fifo_15_tready,
    output ap_fifo_oarg_15_full_n,
    input [C_OUTPUT_FIFO_15_WIDTH-1:0] ap_fifo_oarg_15_din,
    input ap_fifo_oarg_15_write,
    //output FIFO to AXI-Stream interface 16
    output m_axis_fifo_16_tlast,
    output m_axis_fifo_16_tvalid,
    output [C_OUTPUT_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tkeep,
    output [C_OUTPUT_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tstrb,
    output [C_OUTPUT_FIFO_16_DMWIDTH-1:0] m_axis_fifo_16_tdata,
    input m_axis_fifo_16_tready,
    output ap_fifo_oarg_16_full_n,
    input [C_OUTPUT_FIFO_16_WIDTH-1:0] ap_fifo_oarg_16_din,
    input ap_fifo_oarg_16_write,
    //output FIFO to AXI-Stream interface 17
    output m_axis_fifo_17_tlast,
    output m_axis_fifo_17_tvalid,
    output [C_OUTPUT_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tkeep,
    output [C_OUTPUT_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tstrb,
    output [C_OUTPUT_FIFO_17_DMWIDTH-1:0] m_axis_fifo_17_tdata,
    input m_axis_fifo_17_tready,
    output ap_fifo_oarg_17_full_n,
    input [C_OUTPUT_FIFO_17_WIDTH-1:0] ap_fifo_oarg_17_din,
    input ap_fifo_oarg_17_write,
    //output FIFO to AXI-Stream interface 18
    output m_axis_fifo_18_tlast,
    output m_axis_fifo_18_tvalid,
    output [C_OUTPUT_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tkeep,
    output [C_OUTPUT_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tstrb,
    output [C_OUTPUT_FIFO_18_DMWIDTH-1:0] m_axis_fifo_18_tdata,
    input m_axis_fifo_18_tready,
    output ap_fifo_oarg_18_full_n,
    input [C_OUTPUT_FIFO_18_WIDTH-1:0] ap_fifo_oarg_18_din,
    input ap_fifo_oarg_18_write,
    //output FIFO to AXI-Stream interface 19
    output m_axis_fifo_19_tlast,
    output m_axis_fifo_19_tvalid,
    output [C_OUTPUT_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tkeep,
    output [C_OUTPUT_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tstrb,
    output [C_OUTPUT_FIFO_19_DMWIDTH-1:0] m_axis_fifo_19_tdata,
    input m_axis_fifo_19_tready,
    output ap_fifo_oarg_19_full_n,
    input [C_OUTPUT_FIFO_19_WIDTH-1:0] ap_fifo_oarg_19_din,
    input ap_fifo_oarg_19_write,
    //output FIFO to AXI-Stream interface 20
    output m_axis_fifo_20_tlast,
    output m_axis_fifo_20_tvalid,
    output [C_OUTPUT_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tkeep,
    output [C_OUTPUT_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tstrb,
    output [C_OUTPUT_FIFO_20_DMWIDTH-1:0] m_axis_fifo_20_tdata,
    input m_axis_fifo_20_tready,
    output ap_fifo_oarg_20_full_n,
    input [C_OUTPUT_FIFO_20_WIDTH-1:0] ap_fifo_oarg_20_din,
    input ap_fifo_oarg_20_write,
    //output FIFO to AXI-Stream interface 21
    output m_axis_fifo_21_tlast,
    output m_axis_fifo_21_tvalid,
    output [C_OUTPUT_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tkeep,
    output [C_OUTPUT_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tstrb,
    output [C_OUTPUT_FIFO_21_DMWIDTH-1:0] m_axis_fifo_21_tdata,
    input m_axis_fifo_21_tready,
    output ap_fifo_oarg_21_full_n,
    input [C_OUTPUT_FIFO_21_WIDTH-1:0] ap_fifo_oarg_21_din,
    input ap_fifo_oarg_21_write,
    //output FIFO to AXI-Stream interface 22
    output m_axis_fifo_22_tlast,
    output m_axis_fifo_22_tvalid,
    output [C_OUTPUT_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tkeep,
    output [C_OUTPUT_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tstrb,
    output [C_OUTPUT_FIFO_22_DMWIDTH-1:0] m_axis_fifo_22_tdata,
    input m_axis_fifo_22_tready,
    output ap_fifo_oarg_22_full_n,
    input [C_OUTPUT_FIFO_22_WIDTH-1:0] ap_fifo_oarg_22_din,
    input ap_fifo_oarg_22_write,
    //output FIFO to AXI-Stream interface 23
    output m_axis_fifo_23_tlast,
    output m_axis_fifo_23_tvalid,
    output [C_OUTPUT_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tkeep,
    output [C_OUTPUT_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tstrb,
    output [C_OUTPUT_FIFO_23_DMWIDTH-1:0] m_axis_fifo_23_tdata,
    input m_axis_fifo_23_tready,
    output ap_fifo_oarg_23_full_n,
    input [C_OUTPUT_FIFO_23_WIDTH-1:0] ap_fifo_oarg_23_din,
    input ap_fifo_oarg_23_write,
    //output FIFO to AXI-Stream interface 24
    output m_axis_fifo_24_tlast,
    output m_axis_fifo_24_tvalid,
    output [C_OUTPUT_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tkeep,
    output [C_OUTPUT_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tstrb,
    output [C_OUTPUT_FIFO_24_DMWIDTH-1:0] m_axis_fifo_24_tdata,
    input m_axis_fifo_24_tready,
    output ap_fifo_oarg_24_full_n,
    input [C_OUTPUT_FIFO_24_WIDTH-1:0] ap_fifo_oarg_24_din,
    input ap_fifo_oarg_24_write,
    //output FIFO to AXI-Stream interface 25
    output m_axis_fifo_25_tlast,
    output m_axis_fifo_25_tvalid,
    output [C_OUTPUT_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tkeep,
    output [C_OUTPUT_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tstrb,
    output [C_OUTPUT_FIFO_25_DMWIDTH-1:0] m_axis_fifo_25_tdata,
    input m_axis_fifo_25_tready,
    output ap_fifo_oarg_25_full_n,
    input [C_OUTPUT_FIFO_25_WIDTH-1:0] ap_fifo_oarg_25_din,
    input ap_fifo_oarg_25_write,
    //output FIFO to AXI-Stream interface 26
    output m_axis_fifo_26_tlast,
    output m_axis_fifo_26_tvalid,
    output [C_OUTPUT_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tkeep,
    output [C_OUTPUT_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tstrb,
    output [C_OUTPUT_FIFO_26_DMWIDTH-1:0] m_axis_fifo_26_tdata,
    input m_axis_fifo_26_tready,
    output ap_fifo_oarg_26_full_n,
    input [C_OUTPUT_FIFO_26_WIDTH-1:0] ap_fifo_oarg_26_din,
    input ap_fifo_oarg_26_write,
    //output FIFO to AXI-Stream interface 27
    output m_axis_fifo_27_tlast,
    output m_axis_fifo_27_tvalid,
    output [C_OUTPUT_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tkeep,
    output [C_OUTPUT_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tstrb,
    output [C_OUTPUT_FIFO_27_DMWIDTH-1:0] m_axis_fifo_27_tdata,
    input m_axis_fifo_27_tready,
    output ap_fifo_oarg_27_full_n,
    input [C_OUTPUT_FIFO_27_WIDTH-1:0] ap_fifo_oarg_27_din,
    input ap_fifo_oarg_27_write,
    //output FIFO to AXI-Stream interface 28
    output m_axis_fifo_28_tlast,
    output m_axis_fifo_28_tvalid,
    output [C_OUTPUT_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tkeep,
    output [C_OUTPUT_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tstrb,
    output [C_OUTPUT_FIFO_28_DMWIDTH-1:0] m_axis_fifo_28_tdata,
    input m_axis_fifo_28_tready,
    output ap_fifo_oarg_28_full_n,
    input [C_OUTPUT_FIFO_28_WIDTH-1:0] ap_fifo_oarg_28_din,
    input ap_fifo_oarg_28_write,
    //output FIFO to AXI-Stream interface 29
    output m_axis_fifo_29_tlast,
    output m_axis_fifo_29_tvalid,
    output [C_OUTPUT_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tkeep,
    output [C_OUTPUT_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tstrb,
    output [C_OUTPUT_FIFO_29_DMWIDTH-1:0] m_axis_fifo_29_tdata,
    input m_axis_fifo_29_tready,
    output ap_fifo_oarg_29_full_n,
    input [C_OUTPUT_FIFO_29_WIDTH-1:0] ap_fifo_oarg_29_din,
    input ap_fifo_oarg_29_write,
    //output FIFO to AXI-Stream interface 30
    output m_axis_fifo_30_tlast,
    output m_axis_fifo_30_tvalid,
    output [C_OUTPUT_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tkeep,
    output [C_OUTPUT_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tstrb,
    output [C_OUTPUT_FIFO_30_DMWIDTH-1:0] m_axis_fifo_30_tdata,
    input m_axis_fifo_30_tready,
    output ap_fifo_oarg_30_full_n,
    input [C_OUTPUT_FIFO_30_WIDTH-1:0] ap_fifo_oarg_30_din,
    input ap_fifo_oarg_30_write,
    //output FIFO to AXI-Stream interface 31
    output m_axis_fifo_31_tlast,
    output m_axis_fifo_31_tvalid,
    output [C_OUTPUT_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tkeep,
    output [C_OUTPUT_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tstrb,
    output [C_OUTPUT_FIFO_31_DMWIDTH-1:0] m_axis_fifo_31_tdata,
    input m_axis_fifo_31_tready,
    output ap_fifo_oarg_31_full_n,
    input [C_OUTPUT_FIFO_31_WIDTH-1:0] ap_fifo_oarg_31_din,
    input ap_fifo_oarg_31_write,
    //output FIFO to AXI-Stream interface 32
    output m_axis_fifo_32_tlast,
    output m_axis_fifo_32_tvalid,
    output [C_OUTPUT_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tkeep,
    output [C_OUTPUT_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tstrb,
    output [C_OUTPUT_FIFO_32_DMWIDTH-1:0] m_axis_fifo_32_tdata,
    input m_axis_fifo_32_tready,
    output ap_fifo_oarg_32_full_n,
    input [C_OUTPUT_FIFO_32_WIDTH-1:0] ap_fifo_oarg_32_din,
    input ap_fifo_oarg_32_write,
    //output FIFO to AXI-Stream interface 33
    output m_axis_fifo_33_tlast,
    output m_axis_fifo_33_tvalid,
    output [C_OUTPUT_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tkeep,
    output [C_OUTPUT_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tstrb,
    output [C_OUTPUT_FIFO_33_DMWIDTH-1:0] m_axis_fifo_33_tdata,
    input m_axis_fifo_33_tready,
    output ap_fifo_oarg_33_full_n,
    input [C_OUTPUT_FIFO_33_WIDTH-1:0] ap_fifo_oarg_33_din,
    input ap_fifo_oarg_33_write,
    //output FIFO to AXI-Stream interface 34
    output m_axis_fifo_34_tlast,
    output m_axis_fifo_34_tvalid,
    output [C_OUTPUT_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tkeep,
    output [C_OUTPUT_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tstrb,
    output [C_OUTPUT_FIFO_34_DMWIDTH-1:0] m_axis_fifo_34_tdata,
    input m_axis_fifo_34_tready,
    output ap_fifo_oarg_34_full_n,
    input [C_OUTPUT_FIFO_34_WIDTH-1:0] ap_fifo_oarg_34_din,
    input ap_fifo_oarg_34_write,
    //output FIFO to AXI-Stream interface 35
    output m_axis_fifo_35_tlast,
    output m_axis_fifo_35_tvalid,
    output [C_OUTPUT_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tkeep,
    output [C_OUTPUT_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tstrb,
    output [C_OUTPUT_FIFO_35_DMWIDTH-1:0] m_axis_fifo_35_tdata,
    input m_axis_fifo_35_tready,
    output ap_fifo_oarg_35_full_n,
    input [C_OUTPUT_FIFO_35_WIDTH-1:0] ap_fifo_oarg_35_din,
    input ap_fifo_oarg_35_write,
    //output FIFO to AXI-Stream interface 36
    output m_axis_fifo_36_tlast,
    output m_axis_fifo_36_tvalid,
    output [C_OUTPUT_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tkeep,
    output [C_OUTPUT_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tstrb,
    output [C_OUTPUT_FIFO_36_DMWIDTH-1:0] m_axis_fifo_36_tdata,
    input m_axis_fifo_36_tready,
    output ap_fifo_oarg_36_full_n,
    input [C_OUTPUT_FIFO_36_WIDTH-1:0] ap_fifo_oarg_36_din,
    input ap_fifo_oarg_36_write,
    //output FIFO to AXI-Stream interface 37
    output m_axis_fifo_37_tlast,
    output m_axis_fifo_37_tvalid,
    output [C_OUTPUT_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tkeep,
    output [C_OUTPUT_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tstrb,
    output [C_OUTPUT_FIFO_37_DMWIDTH-1:0] m_axis_fifo_37_tdata,
    input m_axis_fifo_37_tready,
    output ap_fifo_oarg_37_full_n,
    input [C_OUTPUT_FIFO_37_WIDTH-1:0] ap_fifo_oarg_37_din,
    input ap_fifo_oarg_37_write,
    //output FIFO to AXI-Stream interface 38
    output m_axis_fifo_38_tlast,
    output m_axis_fifo_38_tvalid,
    output [C_OUTPUT_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tkeep,
    output [C_OUTPUT_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tstrb,
    output [C_OUTPUT_FIFO_38_DMWIDTH-1:0] m_axis_fifo_38_tdata,
    input m_axis_fifo_38_tready,
    output ap_fifo_oarg_38_full_n,
    input [C_OUTPUT_FIFO_38_WIDTH-1:0] ap_fifo_oarg_38_din,
    input ap_fifo_oarg_38_write,
    //output FIFO to AXI-Stream interface 39
    output m_axis_fifo_39_tlast,
    output m_axis_fifo_39_tvalid,
    output [C_OUTPUT_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tkeep,
    output [C_OUTPUT_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tstrb,
    output [C_OUTPUT_FIFO_39_DMWIDTH-1:0] m_axis_fifo_39_tdata,
    input m_axis_fifo_39_tready,
    output ap_fifo_oarg_39_full_n,
    input [C_OUTPUT_FIFO_39_WIDTH-1:0] ap_fifo_oarg_39_din,
    input ap_fifo_oarg_39_write,
    //output FIFO to AXI-Stream interface 40
    output m_axis_fifo_40_tlast,
    output m_axis_fifo_40_tvalid,
    output [C_OUTPUT_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tkeep,
    output [C_OUTPUT_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tstrb,
    output [C_OUTPUT_FIFO_40_DMWIDTH-1:0] m_axis_fifo_40_tdata,
    input m_axis_fifo_40_tready,
    output ap_fifo_oarg_40_full_n,
    input [C_OUTPUT_FIFO_40_WIDTH-1:0] ap_fifo_oarg_40_din,
    input ap_fifo_oarg_40_write,
    //output FIFO to AXI-Stream interface 41
    output m_axis_fifo_41_tlast,
    output m_axis_fifo_41_tvalid,
    output [C_OUTPUT_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tkeep,
    output [C_OUTPUT_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tstrb,
    output [C_OUTPUT_FIFO_41_DMWIDTH-1:0] m_axis_fifo_41_tdata,
    input m_axis_fifo_41_tready,
    output ap_fifo_oarg_41_full_n,
    input [C_OUTPUT_FIFO_41_WIDTH-1:0] ap_fifo_oarg_41_din,
    input ap_fifo_oarg_41_write,
    //output FIFO to AXI-Stream interface 42
    output m_axis_fifo_42_tlast,
    output m_axis_fifo_42_tvalid,
    output [C_OUTPUT_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tkeep,
    output [C_OUTPUT_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tstrb,
    output [C_OUTPUT_FIFO_42_DMWIDTH-1:0] m_axis_fifo_42_tdata,
    input m_axis_fifo_42_tready,
    output ap_fifo_oarg_42_full_n,
    input [C_OUTPUT_FIFO_42_WIDTH-1:0] ap_fifo_oarg_42_din,
    input ap_fifo_oarg_42_write,
    //output FIFO to AXI-Stream interface 43
    output m_axis_fifo_43_tlast,
    output m_axis_fifo_43_tvalid,
    output [C_OUTPUT_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tkeep,
    output [C_OUTPUT_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tstrb,
    output [C_OUTPUT_FIFO_43_DMWIDTH-1:0] m_axis_fifo_43_tdata,
    input m_axis_fifo_43_tready,
    output ap_fifo_oarg_43_full_n,
    input [C_OUTPUT_FIFO_43_WIDTH-1:0] ap_fifo_oarg_43_din,
    input ap_fifo_oarg_43_write,
    //output FIFO to AXI-Stream interface 44
    output m_axis_fifo_44_tlast,
    output m_axis_fifo_44_tvalid,
    output [C_OUTPUT_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tkeep,
    output [C_OUTPUT_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tstrb,
    output [C_OUTPUT_FIFO_44_DMWIDTH-1:0] m_axis_fifo_44_tdata,
    input m_axis_fifo_44_tready,
    output ap_fifo_oarg_44_full_n,
    input [C_OUTPUT_FIFO_44_WIDTH-1:0] ap_fifo_oarg_44_din,
    input ap_fifo_oarg_44_write,
    //output FIFO to AXI-Stream interface 45
    output m_axis_fifo_45_tlast,
    output m_axis_fifo_45_tvalid,
    output [C_OUTPUT_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tkeep,
    output [C_OUTPUT_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tstrb,
    output [C_OUTPUT_FIFO_45_DMWIDTH-1:0] m_axis_fifo_45_tdata,
    input m_axis_fifo_45_tready,
    output ap_fifo_oarg_45_full_n,
    input [C_OUTPUT_FIFO_45_WIDTH-1:0] ap_fifo_oarg_45_din,
    input ap_fifo_oarg_45_write,
    //output FIFO to AXI-Stream interface 46
    output m_axis_fifo_46_tlast,
    output m_axis_fifo_46_tvalid,
    output [C_OUTPUT_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tkeep,
    output [C_OUTPUT_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tstrb,
    output [C_OUTPUT_FIFO_46_DMWIDTH-1:0] m_axis_fifo_46_tdata,
    input m_axis_fifo_46_tready,
    output ap_fifo_oarg_46_full_n,
    input [C_OUTPUT_FIFO_46_WIDTH-1:0] ap_fifo_oarg_46_din,
    input ap_fifo_oarg_46_write,
    //output FIFO to AXI-Stream interface 47
    output m_axis_fifo_47_tlast,
    output m_axis_fifo_47_tvalid,
    output [C_OUTPUT_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tkeep,
    output [C_OUTPUT_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tstrb,
    output [C_OUTPUT_FIFO_47_DMWIDTH-1:0] m_axis_fifo_47_tdata,
    input m_axis_fifo_47_tready,
    output ap_fifo_oarg_47_full_n,
    input [C_OUTPUT_FIFO_47_WIDTH-1:0] ap_fifo_oarg_47_din,
    input ap_fifo_oarg_47_write,
    //output FIFO to AXI-Stream interface 48
    output m_axis_fifo_48_tlast,
    output m_axis_fifo_48_tvalid,
    output [C_OUTPUT_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tkeep,
    output [C_OUTPUT_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tstrb,
    output [C_OUTPUT_FIFO_48_DMWIDTH-1:0] m_axis_fifo_48_tdata,
    input m_axis_fifo_48_tready,
    output ap_fifo_oarg_48_full_n,
    input [C_OUTPUT_FIFO_48_WIDTH-1:0] ap_fifo_oarg_48_din,
    input ap_fifo_oarg_48_write,
    //output FIFO to AXI-Stream interface 49
    output m_axis_fifo_49_tlast,
    output m_axis_fifo_49_tvalid,
    output [C_OUTPUT_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tkeep,
    output [C_OUTPUT_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tstrb,
    output [C_OUTPUT_FIFO_49_DMWIDTH-1:0] m_axis_fifo_49_tdata,
    input m_axis_fifo_49_tready,
    output ap_fifo_oarg_49_full_n,
    input [C_OUTPUT_FIFO_49_WIDTH-1:0] ap_fifo_oarg_49_din,
    input ap_fifo_oarg_49_write,
    //output FIFO to AXI-Stream interface 50
    output m_axis_fifo_50_tlast,
    output m_axis_fifo_50_tvalid,
    output [C_OUTPUT_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tkeep,
    output [C_OUTPUT_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tstrb,
    output [C_OUTPUT_FIFO_50_DMWIDTH-1:0] m_axis_fifo_50_tdata,
    input m_axis_fifo_50_tready,
    output ap_fifo_oarg_50_full_n,
    input [C_OUTPUT_FIFO_50_WIDTH-1:0] ap_fifo_oarg_50_din,
    input ap_fifo_oarg_50_write,
    //output FIFO to AXI-Stream interface 51
    output m_axis_fifo_51_tlast,
    output m_axis_fifo_51_tvalid,
    output [C_OUTPUT_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tkeep,
    output [C_OUTPUT_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tstrb,
    output [C_OUTPUT_FIFO_51_DMWIDTH-1:0] m_axis_fifo_51_tdata,
    input m_axis_fifo_51_tready,
    output ap_fifo_oarg_51_full_n,
    input [C_OUTPUT_FIFO_51_WIDTH-1:0] ap_fifo_oarg_51_din,
    input ap_fifo_oarg_51_write,
    //output FIFO to AXI-Stream interface 52
    output m_axis_fifo_52_tlast,
    output m_axis_fifo_52_tvalid,
    output [C_OUTPUT_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tkeep,
    output [C_OUTPUT_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tstrb,
    output [C_OUTPUT_FIFO_52_DMWIDTH-1:0] m_axis_fifo_52_tdata,
    input m_axis_fifo_52_tready,
    output ap_fifo_oarg_52_full_n,
    input [C_OUTPUT_FIFO_52_WIDTH-1:0] ap_fifo_oarg_52_din,
    input ap_fifo_oarg_52_write,
    //output FIFO to AXI-Stream interface 53
    output m_axis_fifo_53_tlast,
    output m_axis_fifo_53_tvalid,
    output [C_OUTPUT_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tkeep,
    output [C_OUTPUT_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tstrb,
    output [C_OUTPUT_FIFO_53_DMWIDTH-1:0] m_axis_fifo_53_tdata,
    input m_axis_fifo_53_tready,
    output ap_fifo_oarg_53_full_n,
    input [C_OUTPUT_FIFO_53_WIDTH-1:0] ap_fifo_oarg_53_din,
    input ap_fifo_oarg_53_write,
    //output FIFO to AXI-Stream interface 54
    output m_axis_fifo_54_tlast,
    output m_axis_fifo_54_tvalid,
    output [C_OUTPUT_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tkeep,
    output [C_OUTPUT_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tstrb,
    output [C_OUTPUT_FIFO_54_DMWIDTH-1:0] m_axis_fifo_54_tdata,
    input m_axis_fifo_54_tready,
    output ap_fifo_oarg_54_full_n,
    input [C_OUTPUT_FIFO_54_WIDTH-1:0] ap_fifo_oarg_54_din,
    input ap_fifo_oarg_54_write,
    //output FIFO to AXI-Stream interface 55
    output m_axis_fifo_55_tlast,
    output m_axis_fifo_55_tvalid,
    output [C_OUTPUT_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tkeep,
    output [C_OUTPUT_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tstrb,
    output [C_OUTPUT_FIFO_55_DMWIDTH-1:0] m_axis_fifo_55_tdata,
    input m_axis_fifo_55_tready,
    output ap_fifo_oarg_55_full_n,
    input [C_OUTPUT_FIFO_55_WIDTH-1:0] ap_fifo_oarg_55_din,
    input ap_fifo_oarg_55_write,
    //output FIFO to AXI-Stream interface 56
    output m_axis_fifo_56_tlast,
    output m_axis_fifo_56_tvalid,
    output [C_OUTPUT_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tkeep,
    output [C_OUTPUT_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tstrb,
    output [C_OUTPUT_FIFO_56_DMWIDTH-1:0] m_axis_fifo_56_tdata,
    input m_axis_fifo_56_tready,
    output ap_fifo_oarg_56_full_n,
    input [C_OUTPUT_FIFO_56_WIDTH-1:0] ap_fifo_oarg_56_din,
    input ap_fifo_oarg_56_write,
    //output FIFO to AXI-Stream interface 57
    output m_axis_fifo_57_tlast,
    output m_axis_fifo_57_tvalid,
    output [C_OUTPUT_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tkeep,
    output [C_OUTPUT_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tstrb,
    output [C_OUTPUT_FIFO_57_DMWIDTH-1:0] m_axis_fifo_57_tdata,
    input m_axis_fifo_57_tready,
    output ap_fifo_oarg_57_full_n,
    input [C_OUTPUT_FIFO_57_WIDTH-1:0] ap_fifo_oarg_57_din,
    input ap_fifo_oarg_57_write,
    //output FIFO to AXI-Stream interface 58
    output m_axis_fifo_58_tlast,
    output m_axis_fifo_58_tvalid,
    output [C_OUTPUT_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tkeep,
    output [C_OUTPUT_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tstrb,
    output [C_OUTPUT_FIFO_58_DMWIDTH-1:0] m_axis_fifo_58_tdata,
    input m_axis_fifo_58_tready,
    output ap_fifo_oarg_58_full_n,
    input [C_OUTPUT_FIFO_58_WIDTH-1:0] ap_fifo_oarg_58_din,
    input ap_fifo_oarg_58_write,
    //output FIFO to AXI-Stream interface 59
    output m_axis_fifo_59_tlast,
    output m_axis_fifo_59_tvalid,
    output [C_OUTPUT_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tkeep,
    output [C_OUTPUT_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tstrb,
    output [C_OUTPUT_FIFO_59_DMWIDTH-1:0] m_axis_fifo_59_tdata,
    input m_axis_fifo_59_tready,
    output ap_fifo_oarg_59_full_n,
    input [C_OUTPUT_FIFO_59_WIDTH-1:0] ap_fifo_oarg_59_din,
    input ap_fifo_oarg_59_write,
    //output FIFO to AXI-Stream interface 60
    output m_axis_fifo_60_tlast,
    output m_axis_fifo_60_tvalid,
    output [C_OUTPUT_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tkeep,
    output [C_OUTPUT_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tstrb,
    output [C_OUTPUT_FIFO_60_DMWIDTH-1:0] m_axis_fifo_60_tdata,
    input m_axis_fifo_60_tready,
    output ap_fifo_oarg_60_full_n,
    input [C_OUTPUT_FIFO_60_WIDTH-1:0] ap_fifo_oarg_60_din,
    input ap_fifo_oarg_60_write,
    //output FIFO to AXI-Stream interface 61
    output m_axis_fifo_61_tlast,
    output m_axis_fifo_61_tvalid,
    output [C_OUTPUT_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tkeep,
    output [C_OUTPUT_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tstrb,
    output [C_OUTPUT_FIFO_61_DMWIDTH-1:0] m_axis_fifo_61_tdata,
    input m_axis_fifo_61_tready,
    output ap_fifo_oarg_61_full_n,
    input [C_OUTPUT_FIFO_61_WIDTH-1:0] ap_fifo_oarg_61_din,
    input ap_fifo_oarg_61_write,
    //output FIFO to AXI-Stream interface 62
    output m_axis_fifo_62_tlast,
    output m_axis_fifo_62_tvalid,
    output [C_OUTPUT_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tkeep,
    output [C_OUTPUT_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tstrb,
    output [C_OUTPUT_FIFO_62_DMWIDTH-1:0] m_axis_fifo_62_tdata,
    input m_axis_fifo_62_tready,
    output ap_fifo_oarg_62_full_n,
    input [C_OUTPUT_FIFO_62_WIDTH-1:0] ap_fifo_oarg_62_din,
    input ap_fifo_oarg_62_write,
    //output FIFO to AXI-Stream interface 63
    output m_axis_fifo_63_tlast,
    output m_axis_fifo_63_tvalid,
    output [C_OUTPUT_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tkeep,
    output [C_OUTPUT_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tstrb,
    output [C_OUTPUT_FIFO_63_DMWIDTH-1:0] m_axis_fifo_63_tdata,
    input m_axis_fifo_63_tready,
    output ap_fifo_oarg_63_full_n,
    input [C_OUTPUT_FIFO_63_WIDTH-1:0] ap_fifo_oarg_63_din,
    input ap_fifo_oarg_63_write,
    //output FIFO to AXI-Stream interface 64
    output m_axis_fifo_64_tlast,
    output m_axis_fifo_64_tvalid,
    output [C_OUTPUT_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tkeep,
    output [C_OUTPUT_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tstrb,
    output [C_OUTPUT_FIFO_64_DMWIDTH-1:0] m_axis_fifo_64_tdata,
    input m_axis_fifo_64_tready,
    output ap_fifo_oarg_64_full_n,
    input [C_OUTPUT_FIFO_64_WIDTH-1:0] ap_fifo_oarg_64_din,
    input ap_fifo_oarg_64_write,
    //output FIFO to AXI-Stream interface 65
    output m_axis_fifo_65_tlast,
    output m_axis_fifo_65_tvalid,
    output [C_OUTPUT_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tkeep,
    output [C_OUTPUT_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tstrb,
    output [C_OUTPUT_FIFO_65_DMWIDTH-1:0] m_axis_fifo_65_tdata,
    input m_axis_fifo_65_tready,
    output ap_fifo_oarg_65_full_n,
    input [C_OUTPUT_FIFO_65_WIDTH-1:0] ap_fifo_oarg_65_din,
    input ap_fifo_oarg_65_write,
    //output FIFO to AXI-Stream interface 66
    output m_axis_fifo_66_tlast,
    output m_axis_fifo_66_tvalid,
    output [C_OUTPUT_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tkeep,
    output [C_OUTPUT_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tstrb,
    output [C_OUTPUT_FIFO_66_DMWIDTH-1:0] m_axis_fifo_66_tdata,
    input m_axis_fifo_66_tready,
    output ap_fifo_oarg_66_full_n,
    input [C_OUTPUT_FIFO_66_WIDTH-1:0] ap_fifo_oarg_66_din,
    input ap_fifo_oarg_66_write,
    //output FIFO to AXI-Stream interface 67
    output m_axis_fifo_67_tlast,
    output m_axis_fifo_67_tvalid,
    output [C_OUTPUT_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tkeep,
    output [C_OUTPUT_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tstrb,
    output [C_OUTPUT_FIFO_67_DMWIDTH-1:0] m_axis_fifo_67_tdata,
    input m_axis_fifo_67_tready,
    output ap_fifo_oarg_67_full_n,
    input [C_OUTPUT_FIFO_67_WIDTH-1:0] ap_fifo_oarg_67_din,
    input ap_fifo_oarg_67_write,
    //output FIFO to AXI-Stream interface 68
    output m_axis_fifo_68_tlast,
    output m_axis_fifo_68_tvalid,
    output [C_OUTPUT_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tkeep,
    output [C_OUTPUT_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tstrb,
    output [C_OUTPUT_FIFO_68_DMWIDTH-1:0] m_axis_fifo_68_tdata,
    input m_axis_fifo_68_tready,
    output ap_fifo_oarg_68_full_n,
    input [C_OUTPUT_FIFO_68_WIDTH-1:0] ap_fifo_oarg_68_din,
    input ap_fifo_oarg_68_write,
    //output FIFO to AXI-Stream interface 69
    output m_axis_fifo_69_tlast,
    output m_axis_fifo_69_tvalid,
    output [C_OUTPUT_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tkeep,
    output [C_OUTPUT_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tstrb,
    output [C_OUTPUT_FIFO_69_DMWIDTH-1:0] m_axis_fifo_69_tdata,
    input m_axis_fifo_69_tready,
    output ap_fifo_oarg_69_full_n,
    input [C_OUTPUT_FIFO_69_WIDTH-1:0] ap_fifo_oarg_69_din,
    input ap_fifo_oarg_69_write,
    //output FIFO to AXI-Stream interface 70
    output m_axis_fifo_70_tlast,
    output m_axis_fifo_70_tvalid,
    output [C_OUTPUT_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tkeep,
    output [C_OUTPUT_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tstrb,
    output [C_OUTPUT_FIFO_70_DMWIDTH-1:0] m_axis_fifo_70_tdata,
    input m_axis_fifo_70_tready,
    output ap_fifo_oarg_70_full_n,
    input [C_OUTPUT_FIFO_70_WIDTH-1:0] ap_fifo_oarg_70_din,
    input ap_fifo_oarg_70_write,
    //output FIFO to AXI-Stream interface 71
    output m_axis_fifo_71_tlast,
    output m_axis_fifo_71_tvalid,
    output [C_OUTPUT_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tkeep,
    output [C_OUTPUT_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tstrb,
    output [C_OUTPUT_FIFO_71_DMWIDTH-1:0] m_axis_fifo_71_tdata,
    input m_axis_fifo_71_tready,
    output ap_fifo_oarg_71_full_n,
    input [C_OUTPUT_FIFO_71_WIDTH-1:0] ap_fifo_oarg_71_din,
    input ap_fifo_oarg_71_write,
    //output FIFO to AXI-Stream interface 72
    output m_axis_fifo_72_tlast,
    output m_axis_fifo_72_tvalid,
    output [C_OUTPUT_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tkeep,
    output [C_OUTPUT_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tstrb,
    output [C_OUTPUT_FIFO_72_DMWIDTH-1:0] m_axis_fifo_72_tdata,
    input m_axis_fifo_72_tready,
    output ap_fifo_oarg_72_full_n,
    input [C_OUTPUT_FIFO_72_WIDTH-1:0] ap_fifo_oarg_72_din,
    input ap_fifo_oarg_72_write,
    //output FIFO to AXI-Stream interface 73
    output m_axis_fifo_73_tlast,
    output m_axis_fifo_73_tvalid,
    output [C_OUTPUT_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tkeep,
    output [C_OUTPUT_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tstrb,
    output [C_OUTPUT_FIFO_73_DMWIDTH-1:0] m_axis_fifo_73_tdata,
    input m_axis_fifo_73_tready,
    output ap_fifo_oarg_73_full_n,
    input [C_OUTPUT_FIFO_73_WIDTH-1:0] ap_fifo_oarg_73_din,
    input ap_fifo_oarg_73_write,
    //output FIFO to AXI-Stream interface 74
    output m_axis_fifo_74_tlast,
    output m_axis_fifo_74_tvalid,
    output [C_OUTPUT_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tkeep,
    output [C_OUTPUT_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tstrb,
    output [C_OUTPUT_FIFO_74_DMWIDTH-1:0] m_axis_fifo_74_tdata,
    input m_axis_fifo_74_tready,
    output ap_fifo_oarg_74_full_n,
    input [C_OUTPUT_FIFO_74_WIDTH-1:0] ap_fifo_oarg_74_din,
    input ap_fifo_oarg_74_write,
    //output FIFO to AXI-Stream interface 75
    output m_axis_fifo_75_tlast,
    output m_axis_fifo_75_tvalid,
    output [C_OUTPUT_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tkeep,
    output [C_OUTPUT_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tstrb,
    output [C_OUTPUT_FIFO_75_DMWIDTH-1:0] m_axis_fifo_75_tdata,
    input m_axis_fifo_75_tready,
    output ap_fifo_oarg_75_full_n,
    input [C_OUTPUT_FIFO_75_WIDTH-1:0] ap_fifo_oarg_75_din,
    input ap_fifo_oarg_75_write,
    //output FIFO to AXI-Stream interface 76
    output m_axis_fifo_76_tlast,
    output m_axis_fifo_76_tvalid,
    output [C_OUTPUT_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tkeep,
    output [C_OUTPUT_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tstrb,
    output [C_OUTPUT_FIFO_76_DMWIDTH-1:0] m_axis_fifo_76_tdata,
    input m_axis_fifo_76_tready,
    output ap_fifo_oarg_76_full_n,
    input [C_OUTPUT_FIFO_76_WIDTH-1:0] ap_fifo_oarg_76_din,
    input ap_fifo_oarg_76_write,
    //output FIFO to AXI-Stream interface 77
    output m_axis_fifo_77_tlast,
    output m_axis_fifo_77_tvalid,
    output [C_OUTPUT_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tkeep,
    output [C_OUTPUT_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tstrb,
    output [C_OUTPUT_FIFO_77_DMWIDTH-1:0] m_axis_fifo_77_tdata,
    input m_axis_fifo_77_tready,
    output ap_fifo_oarg_77_full_n,
    input [C_OUTPUT_FIFO_77_WIDTH-1:0] ap_fifo_oarg_77_din,
    input ap_fifo_oarg_77_write,
    //output FIFO to AXI-Stream interface 78
    output m_axis_fifo_78_tlast,
    output m_axis_fifo_78_tvalid,
    output [C_OUTPUT_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tkeep,
    output [C_OUTPUT_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tstrb,
    output [C_OUTPUT_FIFO_78_DMWIDTH-1:0] m_axis_fifo_78_tdata,
    input m_axis_fifo_78_tready,
    output ap_fifo_oarg_78_full_n,
    input [C_OUTPUT_FIFO_78_WIDTH-1:0] ap_fifo_oarg_78_din,
    input ap_fifo_oarg_78_write,
    //output FIFO to AXI-Stream interface 79
    output m_axis_fifo_79_tlast,
    output m_axis_fifo_79_tvalid,
    output [C_OUTPUT_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tkeep,
    output [C_OUTPUT_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tstrb,
    output [C_OUTPUT_FIFO_79_DMWIDTH-1:0] m_axis_fifo_79_tdata,
    input m_axis_fifo_79_tready,
    output ap_fifo_oarg_79_full_n,
    input [C_OUTPUT_FIFO_79_WIDTH-1:0] ap_fifo_oarg_79_din,
    input ap_fifo_oarg_79_write,
    //output FIFO to AXI-Stream interface 80
    output m_axis_fifo_80_tlast,
    output m_axis_fifo_80_tvalid,
    output [C_OUTPUT_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tkeep,
    output [C_OUTPUT_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tstrb,
    output [C_OUTPUT_FIFO_80_DMWIDTH-1:0] m_axis_fifo_80_tdata,
    input m_axis_fifo_80_tready,
    output ap_fifo_oarg_80_full_n,
    input [C_OUTPUT_FIFO_80_WIDTH-1:0] ap_fifo_oarg_80_din,
    input ap_fifo_oarg_80_write,
    //output FIFO to AXI-Stream interface 81
    output m_axis_fifo_81_tlast,
    output m_axis_fifo_81_tvalid,
    output [C_OUTPUT_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tkeep,
    output [C_OUTPUT_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tstrb,
    output [C_OUTPUT_FIFO_81_DMWIDTH-1:0] m_axis_fifo_81_tdata,
    input m_axis_fifo_81_tready,
    output ap_fifo_oarg_81_full_n,
    input [C_OUTPUT_FIFO_81_WIDTH-1:0] ap_fifo_oarg_81_din,
    input ap_fifo_oarg_81_write,
    //output FIFO to AXI-Stream interface 82
    output m_axis_fifo_82_tlast,
    output m_axis_fifo_82_tvalid,
    output [C_OUTPUT_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tkeep,
    output [C_OUTPUT_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tstrb,
    output [C_OUTPUT_FIFO_82_DMWIDTH-1:0] m_axis_fifo_82_tdata,
    input m_axis_fifo_82_tready,
    output ap_fifo_oarg_82_full_n,
    input [C_OUTPUT_FIFO_82_WIDTH-1:0] ap_fifo_oarg_82_din,
    input ap_fifo_oarg_82_write,
    //output FIFO to AXI-Stream interface 83
    output m_axis_fifo_83_tlast,
    output m_axis_fifo_83_tvalid,
    output [C_OUTPUT_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tkeep,
    output [C_OUTPUT_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tstrb,
    output [C_OUTPUT_FIFO_83_DMWIDTH-1:0] m_axis_fifo_83_tdata,
    input m_axis_fifo_83_tready,
    output ap_fifo_oarg_83_full_n,
    input [C_OUTPUT_FIFO_83_WIDTH-1:0] ap_fifo_oarg_83_din,
    input ap_fifo_oarg_83_write,
    //output FIFO to AXI-Stream interface 84
    output m_axis_fifo_84_tlast,
    output m_axis_fifo_84_tvalid,
    output [C_OUTPUT_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tkeep,
    output [C_OUTPUT_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tstrb,
    output [C_OUTPUT_FIFO_84_DMWIDTH-1:0] m_axis_fifo_84_tdata,
    input m_axis_fifo_84_tready,
    output ap_fifo_oarg_84_full_n,
    input [C_OUTPUT_FIFO_84_WIDTH-1:0] ap_fifo_oarg_84_din,
    input ap_fifo_oarg_84_write,
    //output FIFO to AXI-Stream interface 85
    output m_axis_fifo_85_tlast,
    output m_axis_fifo_85_tvalid,
    output [C_OUTPUT_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tkeep,
    output [C_OUTPUT_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tstrb,
    output [C_OUTPUT_FIFO_85_DMWIDTH-1:0] m_axis_fifo_85_tdata,
    input m_axis_fifo_85_tready,
    output ap_fifo_oarg_85_full_n,
    input [C_OUTPUT_FIFO_85_WIDTH-1:0] ap_fifo_oarg_85_din,
    input ap_fifo_oarg_85_write,
    //output FIFO to AXI-Stream interface 86
    output m_axis_fifo_86_tlast,
    output m_axis_fifo_86_tvalid,
    output [C_OUTPUT_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tkeep,
    output [C_OUTPUT_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tstrb,
    output [C_OUTPUT_FIFO_86_DMWIDTH-1:0] m_axis_fifo_86_tdata,
    input m_axis_fifo_86_tready,
    output ap_fifo_oarg_86_full_n,
    input [C_OUTPUT_FIFO_86_WIDTH-1:0] ap_fifo_oarg_86_din,
    input ap_fifo_oarg_86_write,
    //output FIFO to AXI-Stream interface 87
    output m_axis_fifo_87_tlast,
    output m_axis_fifo_87_tvalid,
    output [C_OUTPUT_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tkeep,
    output [C_OUTPUT_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tstrb,
    output [C_OUTPUT_FIFO_87_DMWIDTH-1:0] m_axis_fifo_87_tdata,
    input m_axis_fifo_87_tready,
    output ap_fifo_oarg_87_full_n,
    input [C_OUTPUT_FIFO_87_WIDTH-1:0] ap_fifo_oarg_87_din,
    input ap_fifo_oarg_87_write,
    //output FIFO to AXI-Stream interface 88
    output m_axis_fifo_88_tlast,
    output m_axis_fifo_88_tvalid,
    output [C_OUTPUT_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tkeep,
    output [C_OUTPUT_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tstrb,
    output [C_OUTPUT_FIFO_88_DMWIDTH-1:0] m_axis_fifo_88_tdata,
    input m_axis_fifo_88_tready,
    output ap_fifo_oarg_88_full_n,
    input [C_OUTPUT_FIFO_88_WIDTH-1:0] ap_fifo_oarg_88_din,
    input ap_fifo_oarg_88_write,
    //output FIFO to AXI-Stream interface 89
    output m_axis_fifo_89_tlast,
    output m_axis_fifo_89_tvalid,
    output [C_OUTPUT_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tkeep,
    output [C_OUTPUT_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tstrb,
    output [C_OUTPUT_FIFO_89_DMWIDTH-1:0] m_axis_fifo_89_tdata,
    input m_axis_fifo_89_tready,
    output ap_fifo_oarg_89_full_n,
    input [C_OUTPUT_FIFO_89_WIDTH-1:0] ap_fifo_oarg_89_din,
    input ap_fifo_oarg_89_write,
    //output FIFO to AXI-Stream interface 90
    output m_axis_fifo_90_tlast,
    output m_axis_fifo_90_tvalid,
    output [C_OUTPUT_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tkeep,
    output [C_OUTPUT_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tstrb,
    output [C_OUTPUT_FIFO_90_DMWIDTH-1:0] m_axis_fifo_90_tdata,
    input m_axis_fifo_90_tready,
    output ap_fifo_oarg_90_full_n,
    input [C_OUTPUT_FIFO_90_WIDTH-1:0] ap_fifo_oarg_90_din,
    input ap_fifo_oarg_90_write,
    //output FIFO to AXI-Stream interface 91
    output m_axis_fifo_91_tlast,
    output m_axis_fifo_91_tvalid,
    output [C_OUTPUT_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tkeep,
    output [C_OUTPUT_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tstrb,
    output [C_OUTPUT_FIFO_91_DMWIDTH-1:0] m_axis_fifo_91_tdata,
    input m_axis_fifo_91_tready,
    output ap_fifo_oarg_91_full_n,
    input [C_OUTPUT_FIFO_91_WIDTH-1:0] ap_fifo_oarg_91_din,
    input ap_fifo_oarg_91_write,
    //output FIFO to AXI-Stream interface 92
    output m_axis_fifo_92_tlast,
    output m_axis_fifo_92_tvalid,
    output [C_OUTPUT_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tkeep,
    output [C_OUTPUT_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tstrb,
    output [C_OUTPUT_FIFO_92_DMWIDTH-1:0] m_axis_fifo_92_tdata,
    input m_axis_fifo_92_tready,
    output ap_fifo_oarg_92_full_n,
    input [C_OUTPUT_FIFO_92_WIDTH-1:0] ap_fifo_oarg_92_din,
    input ap_fifo_oarg_92_write,
    //output FIFO to AXI-Stream interface 93
    output m_axis_fifo_93_tlast,
    output m_axis_fifo_93_tvalid,
    output [C_OUTPUT_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tkeep,
    output [C_OUTPUT_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tstrb,
    output [C_OUTPUT_FIFO_93_DMWIDTH-1:0] m_axis_fifo_93_tdata,
    input m_axis_fifo_93_tready,
    output ap_fifo_oarg_93_full_n,
    input [C_OUTPUT_FIFO_93_WIDTH-1:0] ap_fifo_oarg_93_din,
    input ap_fifo_oarg_93_write,
    //output FIFO to AXI-Stream interface 94
    output m_axis_fifo_94_tlast,
    output m_axis_fifo_94_tvalid,
    output [C_OUTPUT_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tkeep,
    output [C_OUTPUT_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tstrb,
    output [C_OUTPUT_FIFO_94_DMWIDTH-1:0] m_axis_fifo_94_tdata,
    input m_axis_fifo_94_tready,
    output ap_fifo_oarg_94_full_n,
    input [C_OUTPUT_FIFO_94_WIDTH-1:0] ap_fifo_oarg_94_din,
    input ap_fifo_oarg_94_write,
    //output FIFO to AXI-Stream interface 95
    output m_axis_fifo_95_tlast,
    output m_axis_fifo_95_tvalid,
    output [C_OUTPUT_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tkeep,
    output [C_OUTPUT_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tstrb,
    output [C_OUTPUT_FIFO_95_DMWIDTH-1:0] m_axis_fifo_95_tdata,
    input m_axis_fifo_95_tready,
    output ap_fifo_oarg_95_full_n,
    input [C_OUTPUT_FIFO_95_WIDTH-1:0] ap_fifo_oarg_95_din,
    input ap_fifo_oarg_95_write,
    //output FIFO to AXI-Stream interface 96
    output m_axis_fifo_96_tlast,
    output m_axis_fifo_96_tvalid,
    output [C_OUTPUT_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tkeep,
    output [C_OUTPUT_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tstrb,
    output [C_OUTPUT_FIFO_96_DMWIDTH-1:0] m_axis_fifo_96_tdata,
    input m_axis_fifo_96_tready,
    output ap_fifo_oarg_96_full_n,
    input [C_OUTPUT_FIFO_96_WIDTH-1:0] ap_fifo_oarg_96_din,
    input ap_fifo_oarg_96_write,
    //output FIFO to AXI-Stream interface 97
    output m_axis_fifo_97_tlast,
    output m_axis_fifo_97_tvalid,
    output [C_OUTPUT_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tkeep,
    output [C_OUTPUT_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tstrb,
    output [C_OUTPUT_FIFO_97_DMWIDTH-1:0] m_axis_fifo_97_tdata,
    input m_axis_fifo_97_tready,
    output ap_fifo_oarg_97_full_n,
    input [C_OUTPUT_FIFO_97_WIDTH-1:0] ap_fifo_oarg_97_din,
    input ap_fifo_oarg_97_write,
    //output FIFO to AXI-Stream interface 98
    output m_axis_fifo_98_tlast,
    output m_axis_fifo_98_tvalid,
    output [C_OUTPUT_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tkeep,
    output [C_OUTPUT_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tstrb,
    output [C_OUTPUT_FIFO_98_DMWIDTH-1:0] m_axis_fifo_98_tdata,
    input m_axis_fifo_98_tready,
    output ap_fifo_oarg_98_full_n,
    input [C_OUTPUT_FIFO_98_WIDTH-1:0] ap_fifo_oarg_98_din,
    input ap_fifo_oarg_98_write,
    //output FIFO to AXI-Stream interface 99
    output m_axis_fifo_99_tlast,
    output m_axis_fifo_99_tvalid,
    output [C_OUTPUT_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tkeep,
    output [C_OUTPUT_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tstrb,
    output [C_OUTPUT_FIFO_99_DMWIDTH-1:0] m_axis_fifo_99_tdata,
    input m_axis_fifo_99_tready,
    output ap_fifo_oarg_99_full_n,
    input [C_OUTPUT_FIFO_99_WIDTH-1:0] ap_fifo_oarg_99_din,
    input ap_fifo_oarg_99_write,
    //output FIFO to AXI-Stream interface 100
    output m_axis_fifo_100_tlast,
    output m_axis_fifo_100_tvalid,
    output [C_OUTPUT_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tkeep,
    output [C_OUTPUT_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tstrb,
    output [C_OUTPUT_FIFO_100_DMWIDTH-1:0] m_axis_fifo_100_tdata,
    input m_axis_fifo_100_tready,
    output ap_fifo_oarg_100_full_n,
    input [C_OUTPUT_FIFO_100_WIDTH-1:0] ap_fifo_oarg_100_din,
    input ap_fifo_oarg_100_write,
    //output FIFO to AXI-Stream interface 101
    output m_axis_fifo_101_tlast,
    output m_axis_fifo_101_tvalid,
    output [C_OUTPUT_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tkeep,
    output [C_OUTPUT_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tstrb,
    output [C_OUTPUT_FIFO_101_DMWIDTH-1:0] m_axis_fifo_101_tdata,
    input m_axis_fifo_101_tready,
    output ap_fifo_oarg_101_full_n,
    input [C_OUTPUT_FIFO_101_WIDTH-1:0] ap_fifo_oarg_101_din,
    input ap_fifo_oarg_101_write,
    //output FIFO to AXI-Stream interface 102
    output m_axis_fifo_102_tlast,
    output m_axis_fifo_102_tvalid,
    output [C_OUTPUT_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tkeep,
    output [C_OUTPUT_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tstrb,
    output [C_OUTPUT_FIFO_102_DMWIDTH-1:0] m_axis_fifo_102_tdata,
    input m_axis_fifo_102_tready,
    output ap_fifo_oarg_102_full_n,
    input [C_OUTPUT_FIFO_102_WIDTH-1:0] ap_fifo_oarg_102_din,
    input ap_fifo_oarg_102_write,
    //output FIFO to AXI-Stream interface 103
    output m_axis_fifo_103_tlast,
    output m_axis_fifo_103_tvalid,
    output [C_OUTPUT_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tkeep,
    output [C_OUTPUT_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tstrb,
    output [C_OUTPUT_FIFO_103_DMWIDTH-1:0] m_axis_fifo_103_tdata,
    input m_axis_fifo_103_tready,
    output ap_fifo_oarg_103_full_n,
    input [C_OUTPUT_FIFO_103_WIDTH-1:0] ap_fifo_oarg_103_din,
    input ap_fifo_oarg_103_write,
    //output FIFO to AXI-Stream interface 104
    output m_axis_fifo_104_tlast,
    output m_axis_fifo_104_tvalid,
    output [C_OUTPUT_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tkeep,
    output [C_OUTPUT_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tstrb,
    output [C_OUTPUT_FIFO_104_DMWIDTH-1:0] m_axis_fifo_104_tdata,
    input m_axis_fifo_104_tready,
    output ap_fifo_oarg_104_full_n,
    input [C_OUTPUT_FIFO_104_WIDTH-1:0] ap_fifo_oarg_104_din,
    input ap_fifo_oarg_104_write,
    //output FIFO to AXI-Stream interface 105
    output m_axis_fifo_105_tlast,
    output m_axis_fifo_105_tvalid,
    output [C_OUTPUT_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tkeep,
    output [C_OUTPUT_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tstrb,
    output [C_OUTPUT_FIFO_105_DMWIDTH-1:0] m_axis_fifo_105_tdata,
    input m_axis_fifo_105_tready,
    output ap_fifo_oarg_105_full_n,
    input [C_OUTPUT_FIFO_105_WIDTH-1:0] ap_fifo_oarg_105_din,
    input ap_fifo_oarg_105_write,
    //output FIFO to AXI-Stream interface 106
    output m_axis_fifo_106_tlast,
    output m_axis_fifo_106_tvalid,
    output [C_OUTPUT_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tkeep,
    output [C_OUTPUT_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tstrb,
    output [C_OUTPUT_FIFO_106_DMWIDTH-1:0] m_axis_fifo_106_tdata,
    input m_axis_fifo_106_tready,
    output ap_fifo_oarg_106_full_n,
    input [C_OUTPUT_FIFO_106_WIDTH-1:0] ap_fifo_oarg_106_din,
    input ap_fifo_oarg_106_write,
    //output FIFO to AXI-Stream interface 107
    output m_axis_fifo_107_tlast,
    output m_axis_fifo_107_tvalid,
    output [C_OUTPUT_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tkeep,
    output [C_OUTPUT_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tstrb,
    output [C_OUTPUT_FIFO_107_DMWIDTH-1:0] m_axis_fifo_107_tdata,
    input m_axis_fifo_107_tready,
    output ap_fifo_oarg_107_full_n,
    input [C_OUTPUT_FIFO_107_WIDTH-1:0] ap_fifo_oarg_107_din,
    input ap_fifo_oarg_107_write,
    //output FIFO to AXI-Stream interface 108
    output m_axis_fifo_108_tlast,
    output m_axis_fifo_108_tvalid,
    output [C_OUTPUT_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tkeep,
    output [C_OUTPUT_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tstrb,
    output [C_OUTPUT_FIFO_108_DMWIDTH-1:0] m_axis_fifo_108_tdata,
    input m_axis_fifo_108_tready,
    output ap_fifo_oarg_108_full_n,
    input [C_OUTPUT_FIFO_108_WIDTH-1:0] ap_fifo_oarg_108_din,
    input ap_fifo_oarg_108_write,
    //output FIFO to AXI-Stream interface 109
    output m_axis_fifo_109_tlast,
    output m_axis_fifo_109_tvalid,
    output [C_OUTPUT_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tkeep,
    output [C_OUTPUT_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tstrb,
    output [C_OUTPUT_FIFO_109_DMWIDTH-1:0] m_axis_fifo_109_tdata,
    input m_axis_fifo_109_tready,
    output ap_fifo_oarg_109_full_n,
    input [C_OUTPUT_FIFO_109_WIDTH-1:0] ap_fifo_oarg_109_din,
    input ap_fifo_oarg_109_write,
    //output FIFO to AXI-Stream interface 110
    output m_axis_fifo_110_tlast,
    output m_axis_fifo_110_tvalid,
    output [C_OUTPUT_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tkeep,
    output [C_OUTPUT_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tstrb,
    output [C_OUTPUT_FIFO_110_DMWIDTH-1:0] m_axis_fifo_110_tdata,
    input m_axis_fifo_110_tready,
    output ap_fifo_oarg_110_full_n,
    input [C_OUTPUT_FIFO_110_WIDTH-1:0] ap_fifo_oarg_110_din,
    input ap_fifo_oarg_110_write,
    //output FIFO to AXI-Stream interface 111
    output m_axis_fifo_111_tlast,
    output m_axis_fifo_111_tvalid,
    output [C_OUTPUT_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tkeep,
    output [C_OUTPUT_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tstrb,
    output [C_OUTPUT_FIFO_111_DMWIDTH-1:0] m_axis_fifo_111_tdata,
    input m_axis_fifo_111_tready,
    output ap_fifo_oarg_111_full_n,
    input [C_OUTPUT_FIFO_111_WIDTH-1:0] ap_fifo_oarg_111_din,
    input ap_fifo_oarg_111_write,
    //output FIFO to AXI-Stream interface 112
    output m_axis_fifo_112_tlast,
    output m_axis_fifo_112_tvalid,
    output [C_OUTPUT_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tkeep,
    output [C_OUTPUT_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tstrb,
    output [C_OUTPUT_FIFO_112_DMWIDTH-1:0] m_axis_fifo_112_tdata,
    input m_axis_fifo_112_tready,
    output ap_fifo_oarg_112_full_n,
    input [C_OUTPUT_FIFO_112_WIDTH-1:0] ap_fifo_oarg_112_din,
    input ap_fifo_oarg_112_write,
    //output FIFO to AXI-Stream interface 113
    output m_axis_fifo_113_tlast,
    output m_axis_fifo_113_tvalid,
    output [C_OUTPUT_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tkeep,
    output [C_OUTPUT_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tstrb,
    output [C_OUTPUT_FIFO_113_DMWIDTH-1:0] m_axis_fifo_113_tdata,
    input m_axis_fifo_113_tready,
    output ap_fifo_oarg_113_full_n,
    input [C_OUTPUT_FIFO_113_WIDTH-1:0] ap_fifo_oarg_113_din,
    input ap_fifo_oarg_113_write,
    //output FIFO to AXI-Stream interface 114
    output m_axis_fifo_114_tlast,
    output m_axis_fifo_114_tvalid,
    output [C_OUTPUT_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tkeep,
    output [C_OUTPUT_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tstrb,
    output [C_OUTPUT_FIFO_114_DMWIDTH-1:0] m_axis_fifo_114_tdata,
    input m_axis_fifo_114_tready,
    output ap_fifo_oarg_114_full_n,
    input [C_OUTPUT_FIFO_114_WIDTH-1:0] ap_fifo_oarg_114_din,
    input ap_fifo_oarg_114_write,
    //output FIFO to AXI-Stream interface 115
    output m_axis_fifo_115_tlast,
    output m_axis_fifo_115_tvalid,
    output [C_OUTPUT_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tkeep,
    output [C_OUTPUT_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tstrb,
    output [C_OUTPUT_FIFO_115_DMWIDTH-1:0] m_axis_fifo_115_tdata,
    input m_axis_fifo_115_tready,
    output ap_fifo_oarg_115_full_n,
    input [C_OUTPUT_FIFO_115_WIDTH-1:0] ap_fifo_oarg_115_din,
    input ap_fifo_oarg_115_write,
    //output FIFO to AXI-Stream interface 116
    output m_axis_fifo_116_tlast,
    output m_axis_fifo_116_tvalid,
    output [C_OUTPUT_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tkeep,
    output [C_OUTPUT_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tstrb,
    output [C_OUTPUT_FIFO_116_DMWIDTH-1:0] m_axis_fifo_116_tdata,
    input m_axis_fifo_116_tready,
    output ap_fifo_oarg_116_full_n,
    input [C_OUTPUT_FIFO_116_WIDTH-1:0] ap_fifo_oarg_116_din,
    input ap_fifo_oarg_116_write,
    //output FIFO to AXI-Stream interface 117
    output m_axis_fifo_117_tlast,
    output m_axis_fifo_117_tvalid,
    output [C_OUTPUT_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tkeep,
    output [C_OUTPUT_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tstrb,
    output [C_OUTPUT_FIFO_117_DMWIDTH-1:0] m_axis_fifo_117_tdata,
    input m_axis_fifo_117_tready,
    output ap_fifo_oarg_117_full_n,
    input [C_OUTPUT_FIFO_117_WIDTH-1:0] ap_fifo_oarg_117_din,
    input ap_fifo_oarg_117_write,
    //output FIFO to AXI-Stream interface 118
    output m_axis_fifo_118_tlast,
    output m_axis_fifo_118_tvalid,
    output [C_OUTPUT_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tkeep,
    output [C_OUTPUT_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tstrb,
    output [C_OUTPUT_FIFO_118_DMWIDTH-1:0] m_axis_fifo_118_tdata,
    input m_axis_fifo_118_tready,
    output ap_fifo_oarg_118_full_n,
    input [C_OUTPUT_FIFO_118_WIDTH-1:0] ap_fifo_oarg_118_din,
    input ap_fifo_oarg_118_write,
    //output FIFO to AXI-Stream interface 119
    output m_axis_fifo_119_tlast,
    output m_axis_fifo_119_tvalid,
    output [C_OUTPUT_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tkeep,
    output [C_OUTPUT_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tstrb,
    output [C_OUTPUT_FIFO_119_DMWIDTH-1:0] m_axis_fifo_119_tdata,
    input m_axis_fifo_119_tready,
    output ap_fifo_oarg_119_full_n,
    input [C_OUTPUT_FIFO_119_WIDTH-1:0] ap_fifo_oarg_119_din,
    input ap_fifo_oarg_119_write,
    //output FIFO to AXI-Stream interface 120
    output m_axis_fifo_120_tlast,
    output m_axis_fifo_120_tvalid,
    output [C_OUTPUT_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tkeep,
    output [C_OUTPUT_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tstrb,
    output [C_OUTPUT_FIFO_120_DMWIDTH-1:0] m_axis_fifo_120_tdata,
    input m_axis_fifo_120_tready,
    output ap_fifo_oarg_120_full_n,
    input [C_OUTPUT_FIFO_120_WIDTH-1:0] ap_fifo_oarg_120_din,
    input ap_fifo_oarg_120_write,
    //output FIFO to AXI-Stream interface 121
    output m_axis_fifo_121_tlast,
    output m_axis_fifo_121_tvalid,
    output [C_OUTPUT_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tkeep,
    output [C_OUTPUT_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tstrb,
    output [C_OUTPUT_FIFO_121_DMWIDTH-1:0] m_axis_fifo_121_tdata,
    input m_axis_fifo_121_tready,
    output ap_fifo_oarg_121_full_n,
    input [C_OUTPUT_FIFO_121_WIDTH-1:0] ap_fifo_oarg_121_din,
    input ap_fifo_oarg_121_write,
    //output FIFO to AXI-Stream interface 122
    output m_axis_fifo_122_tlast,
    output m_axis_fifo_122_tvalid,
    output [C_OUTPUT_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tkeep,
    output [C_OUTPUT_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tstrb,
    output [C_OUTPUT_FIFO_122_DMWIDTH-1:0] m_axis_fifo_122_tdata,
    input m_axis_fifo_122_tready,
    output ap_fifo_oarg_122_full_n,
    input [C_OUTPUT_FIFO_122_WIDTH-1:0] ap_fifo_oarg_122_din,
    input ap_fifo_oarg_122_write,
    //output FIFO to AXI-Stream interface 123
    output m_axis_fifo_123_tlast,
    output m_axis_fifo_123_tvalid,
    output [C_OUTPUT_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tkeep,
    output [C_OUTPUT_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tstrb,
    output [C_OUTPUT_FIFO_123_DMWIDTH-1:0] m_axis_fifo_123_tdata,
    input m_axis_fifo_123_tready,
    output ap_fifo_oarg_123_full_n,
    input [C_OUTPUT_FIFO_123_WIDTH-1:0] ap_fifo_oarg_123_din,
    input ap_fifo_oarg_123_write,
    //output FIFO to AXI-Stream interface 124
    output m_axis_fifo_124_tlast,
    output m_axis_fifo_124_tvalid,
    output [C_OUTPUT_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tkeep,
    output [C_OUTPUT_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tstrb,
    output [C_OUTPUT_FIFO_124_DMWIDTH-1:0] m_axis_fifo_124_tdata,
    input m_axis_fifo_124_tready,
    output ap_fifo_oarg_124_full_n,
    input [C_OUTPUT_FIFO_124_WIDTH-1:0] ap_fifo_oarg_124_din,
    input ap_fifo_oarg_124_write,
    //output FIFO to AXI-Stream interface 125
    output m_axis_fifo_125_tlast,
    output m_axis_fifo_125_tvalid,
    output [C_OUTPUT_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tkeep,
    output [C_OUTPUT_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tstrb,
    output [C_OUTPUT_FIFO_125_DMWIDTH-1:0] m_axis_fifo_125_tdata,
    input m_axis_fifo_125_tready,
    output ap_fifo_oarg_125_full_n,
    input [C_OUTPUT_FIFO_125_WIDTH-1:0] ap_fifo_oarg_125_din,
    input ap_fifo_oarg_125_write,
    //output FIFO to AXI-Stream interface 126
    output m_axis_fifo_126_tlast,
    output m_axis_fifo_126_tvalid,
    output [C_OUTPUT_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tkeep,
    output [C_OUTPUT_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tstrb,
    output [C_OUTPUT_FIFO_126_DMWIDTH-1:0] m_axis_fifo_126_tdata,
    input m_axis_fifo_126_tready,
    output ap_fifo_oarg_126_full_n,
    input [C_OUTPUT_FIFO_126_WIDTH-1:0] ap_fifo_oarg_126_din,
    input ap_fifo_oarg_126_write,
    //output FIFO to AXI-Stream interface 127
    output m_axis_fifo_127_tlast,
    output m_axis_fifo_127_tvalid,
    output [C_OUTPUT_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tkeep,
    output [C_OUTPUT_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tstrb,
    output [C_OUTPUT_FIFO_127_DMWIDTH-1:0] m_axis_fifo_127_tdata,
    input m_axis_fifo_127_tready,
    output ap_fifo_oarg_127_full_n,
    input [C_OUTPUT_FIFO_127_WIDTH-1:0] ap_fifo_oarg_127_din,
    input ap_fifo_oarg_127_write,
    //-----------------------------------------------------
    //input AXI-Stream to BRAM interface 0
    input s_axis_bram_0_tlast,
    input s_axis_bram_0_tvalid,
    input [C_INPUT_BRAM_0_DMWIDTH/8-1:0] s_axis_bram_0_tkeep,
    input [C_INPUT_BRAM_0_DMWIDTH/8-1:0] s_axis_bram_0_tstrb,
    input [C_INPUT_BRAM_0_DMWIDTH-1:0] s_axis_bram_0_tdata,
    output s_axis_bram_0_tready,
    input [C_INPUT_BRAM_0_ADDR_WIDTH-1:0] ap_bram_iarg_0_addr0,
    input [C_INPUT_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_din0,
    output [C_INPUT_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_dout0,
    input ap_bram_iarg_0_clk0,
    input ap_bram_iarg_0_rst0,
    input [C_INPUT_BRAM_0_WIDTH/8-1:0] ap_bram_iarg_0_we0,
    input ap_bram_iarg_0_en0,
    input [C_INPUT_BRAM_0_ADDR_WIDTH-1:0] ap_bram_iarg_0_addr1,
    input [C_INPUT_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_din1,
    output [C_INPUT_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_dout1,
    input ap_bram_iarg_0_clk1,
    input ap_bram_iarg_0_rst1,
    input [C_INPUT_BRAM_0_WIDTH/8-1:0] ap_bram_iarg_0_we1,
    input ap_bram_iarg_0_en1,
    //input AXI-Stream to BRAM interface 1
    input s_axis_bram_1_tlast,
    input s_axis_bram_1_tvalid,
    input [C_INPUT_BRAM_1_DMWIDTH/8-1:0] s_axis_bram_1_tkeep,
    input [C_INPUT_BRAM_1_DMWIDTH/8-1:0] s_axis_bram_1_tstrb,
    input [C_INPUT_BRAM_1_DMWIDTH-1:0] s_axis_bram_1_tdata,
    output s_axis_bram_1_tready,
    input [C_INPUT_BRAM_1_ADDR_WIDTH-1:0] ap_bram_iarg_1_addr0,
    input [C_INPUT_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_din0,
    output [C_INPUT_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_dout0,
    input ap_bram_iarg_1_clk0,
    input ap_bram_iarg_1_rst0,
    input [C_INPUT_BRAM_1_WIDTH/8-1:0] ap_bram_iarg_1_we0,
    input ap_bram_iarg_1_en0,
    input [C_INPUT_BRAM_1_ADDR_WIDTH-1:0] ap_bram_iarg_1_addr1,
    input [C_INPUT_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_din1,
    output [C_INPUT_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_dout1,
    input ap_bram_iarg_1_clk1,
    input ap_bram_iarg_1_rst1,
    input [C_INPUT_BRAM_1_WIDTH/8-1:0] ap_bram_iarg_1_we1,
    input ap_bram_iarg_1_en1,
    //input AXI-Stream to BRAM interface 2
    input s_axis_bram_2_tlast,
    input s_axis_bram_2_tvalid,
    input [C_INPUT_BRAM_2_DMWIDTH/8-1:0] s_axis_bram_2_tkeep,
    input [C_INPUT_BRAM_2_DMWIDTH/8-1:0] s_axis_bram_2_tstrb,
    input [C_INPUT_BRAM_2_DMWIDTH-1:0] s_axis_bram_2_tdata,
    output s_axis_bram_2_tready,
    input [C_INPUT_BRAM_2_ADDR_WIDTH-1:0] ap_bram_iarg_2_addr0,
    input [C_INPUT_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_din0,
    output [C_INPUT_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_dout0,
    input ap_bram_iarg_2_clk0,
    input ap_bram_iarg_2_rst0,
    input [C_INPUT_BRAM_2_WIDTH/8-1:0] ap_bram_iarg_2_we0,
    input ap_bram_iarg_2_en0,
    input [C_INPUT_BRAM_2_ADDR_WIDTH-1:0] ap_bram_iarg_2_addr1,
    input [C_INPUT_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_din1,
    output [C_INPUT_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_dout1,
    input ap_bram_iarg_2_clk1,
    input ap_bram_iarg_2_rst1,
    input [C_INPUT_BRAM_2_WIDTH/8-1:0] ap_bram_iarg_2_we1,
    input ap_bram_iarg_2_en1,
    //input AXI-Stream to BRAM interface 3
    input s_axis_bram_3_tlast,
    input s_axis_bram_3_tvalid,
    input [C_INPUT_BRAM_3_DMWIDTH/8-1:0] s_axis_bram_3_tkeep,
    input [C_INPUT_BRAM_3_DMWIDTH/8-1:0] s_axis_bram_3_tstrb,
    input [C_INPUT_BRAM_3_DMWIDTH-1:0] s_axis_bram_3_tdata,
    output s_axis_bram_3_tready,
    input [C_INPUT_BRAM_3_ADDR_WIDTH-1:0] ap_bram_iarg_3_addr0,
    input [C_INPUT_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_din0,
    output [C_INPUT_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_dout0,
    input ap_bram_iarg_3_clk0,
    input ap_bram_iarg_3_rst0,
    input [C_INPUT_BRAM_3_WIDTH/8-1:0] ap_bram_iarg_3_we0,
    input ap_bram_iarg_3_en0,
    input [C_INPUT_BRAM_3_ADDR_WIDTH-1:0] ap_bram_iarg_3_addr1,
    input [C_INPUT_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_din1,
    output [C_INPUT_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_dout1,
    input ap_bram_iarg_3_clk1,
    input ap_bram_iarg_3_rst1,
    input [C_INPUT_BRAM_3_WIDTH/8-1:0] ap_bram_iarg_3_we1,
    input ap_bram_iarg_3_en1,
    //input AXI-Stream to BRAM interface 4
    input s_axis_bram_4_tlast,
    input s_axis_bram_4_tvalid,
    input [C_INPUT_BRAM_4_DMWIDTH/8-1:0] s_axis_bram_4_tkeep,
    input [C_INPUT_BRAM_4_DMWIDTH/8-1:0] s_axis_bram_4_tstrb,
    input [C_INPUT_BRAM_4_DMWIDTH-1:0] s_axis_bram_4_tdata,
    output s_axis_bram_4_tready,
    input [C_INPUT_BRAM_4_ADDR_WIDTH-1:0] ap_bram_iarg_4_addr0,
    input [C_INPUT_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_din0,
    output [C_INPUT_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_dout0,
    input ap_bram_iarg_4_clk0,
    input ap_bram_iarg_4_rst0,
    input [C_INPUT_BRAM_4_WIDTH/8-1:0] ap_bram_iarg_4_we0,
    input ap_bram_iarg_4_en0,
    input [C_INPUT_BRAM_4_ADDR_WIDTH-1:0] ap_bram_iarg_4_addr1,
    input [C_INPUT_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_din1,
    output [C_INPUT_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_dout1,
    input ap_bram_iarg_4_clk1,
    input ap_bram_iarg_4_rst1,
    input [C_INPUT_BRAM_4_WIDTH/8-1:0] ap_bram_iarg_4_we1,
    input ap_bram_iarg_4_en1,
    //input AXI-Stream to BRAM interface 5
    input s_axis_bram_5_tlast,
    input s_axis_bram_5_tvalid,
    input [C_INPUT_BRAM_5_DMWIDTH/8-1:0] s_axis_bram_5_tkeep,
    input [C_INPUT_BRAM_5_DMWIDTH/8-1:0] s_axis_bram_5_tstrb,
    input [C_INPUT_BRAM_5_DMWIDTH-1:0] s_axis_bram_5_tdata,
    output s_axis_bram_5_tready,
    input [C_INPUT_BRAM_5_ADDR_WIDTH-1:0] ap_bram_iarg_5_addr0,
    input [C_INPUT_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_din0,
    output [C_INPUT_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_dout0,
    input ap_bram_iarg_5_clk0,
    input ap_bram_iarg_5_rst0,
    input [C_INPUT_BRAM_5_WIDTH/8-1:0] ap_bram_iarg_5_we0,
    input ap_bram_iarg_5_en0,
    input [C_INPUT_BRAM_5_ADDR_WIDTH-1:0] ap_bram_iarg_5_addr1,
    input [C_INPUT_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_din1,
    output [C_INPUT_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_dout1,
    input ap_bram_iarg_5_clk1,
    input ap_bram_iarg_5_rst1,
    input [C_INPUT_BRAM_5_WIDTH/8-1:0] ap_bram_iarg_5_we1,
    input ap_bram_iarg_5_en1,
    //input AXI-Stream to BRAM interface 6
    input s_axis_bram_6_tlast,
    input s_axis_bram_6_tvalid,
    input [C_INPUT_BRAM_6_DMWIDTH/8-1:0] s_axis_bram_6_tkeep,
    input [C_INPUT_BRAM_6_DMWIDTH/8-1:0] s_axis_bram_6_tstrb,
    input [C_INPUT_BRAM_6_DMWIDTH-1:0] s_axis_bram_6_tdata,
    output s_axis_bram_6_tready,
    input [C_INPUT_BRAM_6_ADDR_WIDTH-1:0] ap_bram_iarg_6_addr0,
    input [C_INPUT_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_din0,
    output [C_INPUT_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_dout0,
    input ap_bram_iarg_6_clk0,
    input ap_bram_iarg_6_rst0,
    input [C_INPUT_BRAM_6_WIDTH/8-1:0] ap_bram_iarg_6_we0,
    input ap_bram_iarg_6_en0,
    input [C_INPUT_BRAM_6_ADDR_WIDTH-1:0] ap_bram_iarg_6_addr1,
    input [C_INPUT_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_din1,
    output [C_INPUT_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_dout1,
    input ap_bram_iarg_6_clk1,
    input ap_bram_iarg_6_rst1,
    input [C_INPUT_BRAM_6_WIDTH/8-1:0] ap_bram_iarg_6_we1,
    input ap_bram_iarg_6_en1,
    //input AXI-Stream to BRAM interface 7
    input s_axis_bram_7_tlast,
    input s_axis_bram_7_tvalid,
    input [C_INPUT_BRAM_7_DMWIDTH/8-1:0] s_axis_bram_7_tkeep,
    input [C_INPUT_BRAM_7_DMWIDTH/8-1:0] s_axis_bram_7_tstrb,
    input [C_INPUT_BRAM_7_DMWIDTH-1:0] s_axis_bram_7_tdata,
    output s_axis_bram_7_tready,
    input [C_INPUT_BRAM_7_ADDR_WIDTH-1:0] ap_bram_iarg_7_addr0,
    input [C_INPUT_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_din0,
    output [C_INPUT_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_dout0,
    input ap_bram_iarg_7_clk0,
    input ap_bram_iarg_7_rst0,
    input [C_INPUT_BRAM_7_WIDTH/8-1:0] ap_bram_iarg_7_we0,
    input ap_bram_iarg_7_en0,
    input [C_INPUT_BRAM_7_ADDR_WIDTH-1:0] ap_bram_iarg_7_addr1,
    input [C_INPUT_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_din1,
    output [C_INPUT_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_dout1,
    input ap_bram_iarg_7_clk1,
    input ap_bram_iarg_7_rst1,
    input [C_INPUT_BRAM_7_WIDTH/8-1:0] ap_bram_iarg_7_we1,
    input ap_bram_iarg_7_en1,
    //input AXI-Stream to BRAM interface 8
    input s_axis_bram_8_tlast,
    input s_axis_bram_8_tvalid,
    input [C_INPUT_BRAM_8_DMWIDTH/8-1:0] s_axis_bram_8_tkeep,
    input [C_INPUT_BRAM_8_DMWIDTH/8-1:0] s_axis_bram_8_tstrb,
    input [C_INPUT_BRAM_8_DMWIDTH-1:0] s_axis_bram_8_tdata,
    output s_axis_bram_8_tready,
    input [C_INPUT_BRAM_8_ADDR_WIDTH-1:0] ap_bram_iarg_8_addr0,
    input [C_INPUT_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_din0,
    output [C_INPUT_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_dout0,
    input ap_bram_iarg_8_clk0,
    input ap_bram_iarg_8_rst0,
    input [C_INPUT_BRAM_8_WIDTH/8-1:0] ap_bram_iarg_8_we0,
    input ap_bram_iarg_8_en0,
    input [C_INPUT_BRAM_8_ADDR_WIDTH-1:0] ap_bram_iarg_8_addr1,
    input [C_INPUT_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_din1,
    output [C_INPUT_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_dout1,
    input ap_bram_iarg_8_clk1,
    input ap_bram_iarg_8_rst1,
    input [C_INPUT_BRAM_8_WIDTH/8-1:0] ap_bram_iarg_8_we1,
    input ap_bram_iarg_8_en1,
    //input AXI-Stream to BRAM interface 9
    input s_axis_bram_9_tlast,
    input s_axis_bram_9_tvalid,
    input [C_INPUT_BRAM_9_DMWIDTH/8-1:0] s_axis_bram_9_tkeep,
    input [C_INPUT_BRAM_9_DMWIDTH/8-1:0] s_axis_bram_9_tstrb,
    input [C_INPUT_BRAM_9_DMWIDTH-1:0] s_axis_bram_9_tdata,
    output s_axis_bram_9_tready,
    input [C_INPUT_BRAM_9_ADDR_WIDTH-1:0] ap_bram_iarg_9_addr0,
    input [C_INPUT_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_din0,
    output [C_INPUT_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_dout0,
    input ap_bram_iarg_9_clk0,
    input ap_bram_iarg_9_rst0,
    input [C_INPUT_BRAM_9_WIDTH/8-1:0] ap_bram_iarg_9_we0,
    input ap_bram_iarg_9_en0,
    input [C_INPUT_BRAM_9_ADDR_WIDTH-1:0] ap_bram_iarg_9_addr1,
    input [C_INPUT_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_din1,
    output [C_INPUT_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_dout1,
    input ap_bram_iarg_9_clk1,
    input ap_bram_iarg_9_rst1,
    input [C_INPUT_BRAM_9_WIDTH/8-1:0] ap_bram_iarg_9_we1,
    input ap_bram_iarg_9_en1,
    //input AXI-Stream to BRAM interface 10
    input s_axis_bram_10_tlast,
    input s_axis_bram_10_tvalid,
    input [C_INPUT_BRAM_10_DMWIDTH/8-1:0] s_axis_bram_10_tkeep,
    input [C_INPUT_BRAM_10_DMWIDTH/8-1:0] s_axis_bram_10_tstrb,
    input [C_INPUT_BRAM_10_DMWIDTH-1:0] s_axis_bram_10_tdata,
    output s_axis_bram_10_tready,
    input [C_INPUT_BRAM_10_ADDR_WIDTH-1:0] ap_bram_iarg_10_addr0,
    input [C_INPUT_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_din0,
    output [C_INPUT_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_dout0,
    input ap_bram_iarg_10_clk0,
    input ap_bram_iarg_10_rst0,
    input [C_INPUT_BRAM_10_WIDTH/8-1:0] ap_bram_iarg_10_we0,
    input ap_bram_iarg_10_en0,
    input [C_INPUT_BRAM_10_ADDR_WIDTH-1:0] ap_bram_iarg_10_addr1,
    input [C_INPUT_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_din1,
    output [C_INPUT_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_dout1,
    input ap_bram_iarg_10_clk1,
    input ap_bram_iarg_10_rst1,
    input [C_INPUT_BRAM_10_WIDTH/8-1:0] ap_bram_iarg_10_we1,
    input ap_bram_iarg_10_en1,
    //input AXI-Stream to BRAM interface 11
    input s_axis_bram_11_tlast,
    input s_axis_bram_11_tvalid,
    input [C_INPUT_BRAM_11_DMWIDTH/8-1:0] s_axis_bram_11_tkeep,
    input [C_INPUT_BRAM_11_DMWIDTH/8-1:0] s_axis_bram_11_tstrb,
    input [C_INPUT_BRAM_11_DMWIDTH-1:0] s_axis_bram_11_tdata,
    output s_axis_bram_11_tready,
    input [C_INPUT_BRAM_11_ADDR_WIDTH-1:0] ap_bram_iarg_11_addr0,
    input [C_INPUT_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_din0,
    output [C_INPUT_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_dout0,
    input ap_bram_iarg_11_clk0,
    input ap_bram_iarg_11_rst0,
    input [C_INPUT_BRAM_11_WIDTH/8-1:0] ap_bram_iarg_11_we0,
    input ap_bram_iarg_11_en0,
    input [C_INPUT_BRAM_11_ADDR_WIDTH-1:0] ap_bram_iarg_11_addr1,
    input [C_INPUT_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_din1,
    output [C_INPUT_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_dout1,
    input ap_bram_iarg_11_clk1,
    input ap_bram_iarg_11_rst1,
    input [C_INPUT_BRAM_11_WIDTH/8-1:0] ap_bram_iarg_11_we1,
    input ap_bram_iarg_11_en1,
    //input AXI-Stream to BRAM interface 12
    input s_axis_bram_12_tlast,
    input s_axis_bram_12_tvalid,
    input [C_INPUT_BRAM_12_DMWIDTH/8-1:0] s_axis_bram_12_tkeep,
    input [C_INPUT_BRAM_12_DMWIDTH/8-1:0] s_axis_bram_12_tstrb,
    input [C_INPUT_BRAM_12_DMWIDTH-1:0] s_axis_bram_12_tdata,
    output s_axis_bram_12_tready,
    input [C_INPUT_BRAM_12_ADDR_WIDTH-1:0] ap_bram_iarg_12_addr0,
    input [C_INPUT_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_din0,
    output [C_INPUT_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_dout0,
    input ap_bram_iarg_12_clk0,
    input ap_bram_iarg_12_rst0,
    input [C_INPUT_BRAM_12_WIDTH/8-1:0] ap_bram_iarg_12_we0,
    input ap_bram_iarg_12_en0,
    input [C_INPUT_BRAM_12_ADDR_WIDTH-1:0] ap_bram_iarg_12_addr1,
    input [C_INPUT_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_din1,
    output [C_INPUT_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_dout1,
    input ap_bram_iarg_12_clk1,
    input ap_bram_iarg_12_rst1,
    input [C_INPUT_BRAM_12_WIDTH/8-1:0] ap_bram_iarg_12_we1,
    input ap_bram_iarg_12_en1,
    //input AXI-Stream to BRAM interface 13
    input s_axis_bram_13_tlast,
    input s_axis_bram_13_tvalid,
    input [C_INPUT_BRAM_13_DMWIDTH/8-1:0] s_axis_bram_13_tkeep,
    input [C_INPUT_BRAM_13_DMWIDTH/8-1:0] s_axis_bram_13_tstrb,
    input [C_INPUT_BRAM_13_DMWIDTH-1:0] s_axis_bram_13_tdata,
    output s_axis_bram_13_tready,
    input [C_INPUT_BRAM_13_ADDR_WIDTH-1:0] ap_bram_iarg_13_addr0,
    input [C_INPUT_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_din0,
    output [C_INPUT_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_dout0,
    input ap_bram_iarg_13_clk0,
    input ap_bram_iarg_13_rst0,
    input [C_INPUT_BRAM_13_WIDTH/8-1:0] ap_bram_iarg_13_we0,
    input ap_bram_iarg_13_en0,
    input [C_INPUT_BRAM_13_ADDR_WIDTH-1:0] ap_bram_iarg_13_addr1,
    input [C_INPUT_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_din1,
    output [C_INPUT_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_dout1,
    input ap_bram_iarg_13_clk1,
    input ap_bram_iarg_13_rst1,
    input [C_INPUT_BRAM_13_WIDTH/8-1:0] ap_bram_iarg_13_we1,
    input ap_bram_iarg_13_en1,
    //input AXI-Stream to BRAM interface 14
    input s_axis_bram_14_tlast,
    input s_axis_bram_14_tvalid,
    input [C_INPUT_BRAM_14_DMWIDTH/8-1:0] s_axis_bram_14_tkeep,
    input [C_INPUT_BRAM_14_DMWIDTH/8-1:0] s_axis_bram_14_tstrb,
    input [C_INPUT_BRAM_14_DMWIDTH-1:0] s_axis_bram_14_tdata,
    output s_axis_bram_14_tready,
    input [C_INPUT_BRAM_14_ADDR_WIDTH-1:0] ap_bram_iarg_14_addr0,
    input [C_INPUT_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_din0,
    output [C_INPUT_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_dout0,
    input ap_bram_iarg_14_clk0,
    input ap_bram_iarg_14_rst0,
    input [C_INPUT_BRAM_14_WIDTH/8-1:0] ap_bram_iarg_14_we0,
    input ap_bram_iarg_14_en0,
    input [C_INPUT_BRAM_14_ADDR_WIDTH-1:0] ap_bram_iarg_14_addr1,
    input [C_INPUT_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_din1,
    output [C_INPUT_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_dout1,
    input ap_bram_iarg_14_clk1,
    input ap_bram_iarg_14_rst1,
    input [C_INPUT_BRAM_14_WIDTH/8-1:0] ap_bram_iarg_14_we1,
    input ap_bram_iarg_14_en1,
    //input AXI-Stream to BRAM interface 15
    input s_axis_bram_15_tlast,
    input s_axis_bram_15_tvalid,
    input [C_INPUT_BRAM_15_DMWIDTH/8-1:0] s_axis_bram_15_tkeep,
    input [C_INPUT_BRAM_15_DMWIDTH/8-1:0] s_axis_bram_15_tstrb,
    input [C_INPUT_BRAM_15_DMWIDTH-1:0] s_axis_bram_15_tdata,
    output s_axis_bram_15_tready,
    input [C_INPUT_BRAM_15_ADDR_WIDTH-1:0] ap_bram_iarg_15_addr0,
    input [C_INPUT_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_din0,
    output [C_INPUT_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_dout0,
    input ap_bram_iarg_15_clk0,
    input ap_bram_iarg_15_rst0,
    input [C_INPUT_BRAM_15_WIDTH/8-1:0] ap_bram_iarg_15_we0,
    input ap_bram_iarg_15_en0,
    input [C_INPUT_BRAM_15_ADDR_WIDTH-1:0] ap_bram_iarg_15_addr1,
    input [C_INPUT_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_din1,
    output [C_INPUT_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_dout1,
    input ap_bram_iarg_15_clk1,
    input ap_bram_iarg_15_rst1,
    input [C_INPUT_BRAM_15_WIDTH/8-1:0] ap_bram_iarg_15_we1,
    input ap_bram_iarg_15_en1,
    //input AXI-Stream to BRAM interface 16
    input s_axis_bram_16_tlast,
    input s_axis_bram_16_tvalid,
    input [C_INPUT_BRAM_16_DMWIDTH/8-1:0] s_axis_bram_16_tkeep,
    input [C_INPUT_BRAM_16_DMWIDTH/8-1:0] s_axis_bram_16_tstrb,
    input [C_INPUT_BRAM_16_DMWIDTH-1:0] s_axis_bram_16_tdata,
    output s_axis_bram_16_tready,
    input [C_INPUT_BRAM_16_ADDR_WIDTH-1:0] ap_bram_iarg_16_addr0,
    input [C_INPUT_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_din0,
    output [C_INPUT_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_dout0,
    input ap_bram_iarg_16_clk0,
    input ap_bram_iarg_16_rst0,
    input [C_INPUT_BRAM_16_WIDTH/8-1:0] ap_bram_iarg_16_we0,
    input ap_bram_iarg_16_en0,
    input [C_INPUT_BRAM_16_ADDR_WIDTH-1:0] ap_bram_iarg_16_addr1,
    input [C_INPUT_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_din1,
    output [C_INPUT_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_dout1,
    input ap_bram_iarg_16_clk1,
    input ap_bram_iarg_16_rst1,
    input [C_INPUT_BRAM_16_WIDTH/8-1:0] ap_bram_iarg_16_we1,
    input ap_bram_iarg_16_en1,
    //input AXI-Stream to BRAM interface 17
    input s_axis_bram_17_tlast,
    input s_axis_bram_17_tvalid,
    input [C_INPUT_BRAM_17_DMWIDTH/8-1:0] s_axis_bram_17_tkeep,
    input [C_INPUT_BRAM_17_DMWIDTH/8-1:0] s_axis_bram_17_tstrb,
    input [C_INPUT_BRAM_17_DMWIDTH-1:0] s_axis_bram_17_tdata,
    output s_axis_bram_17_tready,
    input [C_INPUT_BRAM_17_ADDR_WIDTH-1:0] ap_bram_iarg_17_addr0,
    input [C_INPUT_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_din0,
    output [C_INPUT_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_dout0,
    input ap_bram_iarg_17_clk0,
    input ap_bram_iarg_17_rst0,
    input [C_INPUT_BRAM_17_WIDTH/8-1:0] ap_bram_iarg_17_we0,
    input ap_bram_iarg_17_en0,
    input [C_INPUT_BRAM_17_ADDR_WIDTH-1:0] ap_bram_iarg_17_addr1,
    input [C_INPUT_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_din1,
    output [C_INPUT_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_dout1,
    input ap_bram_iarg_17_clk1,
    input ap_bram_iarg_17_rst1,
    input [C_INPUT_BRAM_17_WIDTH/8-1:0] ap_bram_iarg_17_we1,
    input ap_bram_iarg_17_en1,
    //input AXI-Stream to BRAM interface 18
    input s_axis_bram_18_tlast,
    input s_axis_bram_18_tvalid,
    input [C_INPUT_BRAM_18_DMWIDTH/8-1:0] s_axis_bram_18_tkeep,
    input [C_INPUT_BRAM_18_DMWIDTH/8-1:0] s_axis_bram_18_tstrb,
    input [C_INPUT_BRAM_18_DMWIDTH-1:0] s_axis_bram_18_tdata,
    output s_axis_bram_18_tready,
    input [C_INPUT_BRAM_18_ADDR_WIDTH-1:0] ap_bram_iarg_18_addr0,
    input [C_INPUT_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_din0,
    output [C_INPUT_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_dout0,
    input ap_bram_iarg_18_clk0,
    input ap_bram_iarg_18_rst0,
    input [C_INPUT_BRAM_18_WIDTH/8-1:0] ap_bram_iarg_18_we0,
    input ap_bram_iarg_18_en0,
    input [C_INPUT_BRAM_18_ADDR_WIDTH-1:0] ap_bram_iarg_18_addr1,
    input [C_INPUT_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_din1,
    output [C_INPUT_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_dout1,
    input ap_bram_iarg_18_clk1,
    input ap_bram_iarg_18_rst1,
    input [C_INPUT_BRAM_18_WIDTH/8-1:0] ap_bram_iarg_18_we1,
    input ap_bram_iarg_18_en1,
    //input AXI-Stream to BRAM interface 19
    input s_axis_bram_19_tlast,
    input s_axis_bram_19_tvalid,
    input [C_INPUT_BRAM_19_DMWIDTH/8-1:0] s_axis_bram_19_tkeep,
    input [C_INPUT_BRAM_19_DMWIDTH/8-1:0] s_axis_bram_19_tstrb,
    input [C_INPUT_BRAM_19_DMWIDTH-1:0] s_axis_bram_19_tdata,
    output s_axis_bram_19_tready,
    input [C_INPUT_BRAM_19_ADDR_WIDTH-1:0] ap_bram_iarg_19_addr0,
    input [C_INPUT_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_din0,
    output [C_INPUT_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_dout0,
    input ap_bram_iarg_19_clk0,
    input ap_bram_iarg_19_rst0,
    input [C_INPUT_BRAM_19_WIDTH/8-1:0] ap_bram_iarg_19_we0,
    input ap_bram_iarg_19_en0,
    input [C_INPUT_BRAM_19_ADDR_WIDTH-1:0] ap_bram_iarg_19_addr1,
    input [C_INPUT_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_din1,
    output [C_INPUT_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_dout1,
    input ap_bram_iarg_19_clk1,
    input ap_bram_iarg_19_rst1,
    input [C_INPUT_BRAM_19_WIDTH/8-1:0] ap_bram_iarg_19_we1,
    input ap_bram_iarg_19_en1,
    //input AXI-Stream to BRAM interface 20
    input s_axis_bram_20_tlast,
    input s_axis_bram_20_tvalid,
    input [C_INPUT_BRAM_20_DMWIDTH/8-1:0] s_axis_bram_20_tkeep,
    input [C_INPUT_BRAM_20_DMWIDTH/8-1:0] s_axis_bram_20_tstrb,
    input [C_INPUT_BRAM_20_DMWIDTH-1:0] s_axis_bram_20_tdata,
    output s_axis_bram_20_tready,
    input [C_INPUT_BRAM_20_ADDR_WIDTH-1:0] ap_bram_iarg_20_addr0,
    input [C_INPUT_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_din0,
    output [C_INPUT_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_dout0,
    input ap_bram_iarg_20_clk0,
    input ap_bram_iarg_20_rst0,
    input [C_INPUT_BRAM_20_WIDTH/8-1:0] ap_bram_iarg_20_we0,
    input ap_bram_iarg_20_en0,
    input [C_INPUT_BRAM_20_ADDR_WIDTH-1:0] ap_bram_iarg_20_addr1,
    input [C_INPUT_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_din1,
    output [C_INPUT_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_dout1,
    input ap_bram_iarg_20_clk1,
    input ap_bram_iarg_20_rst1,
    input [C_INPUT_BRAM_20_WIDTH/8-1:0] ap_bram_iarg_20_we1,
    input ap_bram_iarg_20_en1,
    //input AXI-Stream to BRAM interface 21
    input s_axis_bram_21_tlast,
    input s_axis_bram_21_tvalid,
    input [C_INPUT_BRAM_21_DMWIDTH/8-1:0] s_axis_bram_21_tkeep,
    input [C_INPUT_BRAM_21_DMWIDTH/8-1:0] s_axis_bram_21_tstrb,
    input [C_INPUT_BRAM_21_DMWIDTH-1:0] s_axis_bram_21_tdata,
    output s_axis_bram_21_tready,
    input [C_INPUT_BRAM_21_ADDR_WIDTH-1:0] ap_bram_iarg_21_addr0,
    input [C_INPUT_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_din0,
    output [C_INPUT_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_dout0,
    input ap_bram_iarg_21_clk0,
    input ap_bram_iarg_21_rst0,
    input [C_INPUT_BRAM_21_WIDTH/8-1:0] ap_bram_iarg_21_we0,
    input ap_bram_iarg_21_en0,
    input [C_INPUT_BRAM_21_ADDR_WIDTH-1:0] ap_bram_iarg_21_addr1,
    input [C_INPUT_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_din1,
    output [C_INPUT_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_dout1,
    input ap_bram_iarg_21_clk1,
    input ap_bram_iarg_21_rst1,
    input [C_INPUT_BRAM_21_WIDTH/8-1:0] ap_bram_iarg_21_we1,
    input ap_bram_iarg_21_en1,
    //input AXI-Stream to BRAM interface 22
    input s_axis_bram_22_tlast,
    input s_axis_bram_22_tvalid,
    input [C_INPUT_BRAM_22_DMWIDTH/8-1:0] s_axis_bram_22_tkeep,
    input [C_INPUT_BRAM_22_DMWIDTH/8-1:0] s_axis_bram_22_tstrb,
    input [C_INPUT_BRAM_22_DMWIDTH-1:0] s_axis_bram_22_tdata,
    output s_axis_bram_22_tready,
    input [C_INPUT_BRAM_22_ADDR_WIDTH-1:0] ap_bram_iarg_22_addr0,
    input [C_INPUT_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_din0,
    output [C_INPUT_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_dout0,
    input ap_bram_iarg_22_clk0,
    input ap_bram_iarg_22_rst0,
    input [C_INPUT_BRAM_22_WIDTH/8-1:0] ap_bram_iarg_22_we0,
    input ap_bram_iarg_22_en0,
    input [C_INPUT_BRAM_22_ADDR_WIDTH-1:0] ap_bram_iarg_22_addr1,
    input [C_INPUT_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_din1,
    output [C_INPUT_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_dout1,
    input ap_bram_iarg_22_clk1,
    input ap_bram_iarg_22_rst1,
    input [C_INPUT_BRAM_22_WIDTH/8-1:0] ap_bram_iarg_22_we1,
    input ap_bram_iarg_22_en1,
    //input AXI-Stream to BRAM interface 23
    input s_axis_bram_23_tlast,
    input s_axis_bram_23_tvalid,
    input [C_INPUT_BRAM_23_DMWIDTH/8-1:0] s_axis_bram_23_tkeep,
    input [C_INPUT_BRAM_23_DMWIDTH/8-1:0] s_axis_bram_23_tstrb,
    input [C_INPUT_BRAM_23_DMWIDTH-1:0] s_axis_bram_23_tdata,
    output s_axis_bram_23_tready,
    input [C_INPUT_BRAM_23_ADDR_WIDTH-1:0] ap_bram_iarg_23_addr0,
    input [C_INPUT_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_din0,
    output [C_INPUT_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_dout0,
    input ap_bram_iarg_23_clk0,
    input ap_bram_iarg_23_rst0,
    input [C_INPUT_BRAM_23_WIDTH/8-1:0] ap_bram_iarg_23_we0,
    input ap_bram_iarg_23_en0,
    input [C_INPUT_BRAM_23_ADDR_WIDTH-1:0] ap_bram_iarg_23_addr1,
    input [C_INPUT_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_din1,
    output [C_INPUT_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_dout1,
    input ap_bram_iarg_23_clk1,
    input ap_bram_iarg_23_rst1,
    input [C_INPUT_BRAM_23_WIDTH/8-1:0] ap_bram_iarg_23_we1,
    input ap_bram_iarg_23_en1,
    //input AXI-Stream to BRAM interface 24
    input s_axis_bram_24_tlast,
    input s_axis_bram_24_tvalid,
    input [C_INPUT_BRAM_24_DMWIDTH/8-1:0] s_axis_bram_24_tkeep,
    input [C_INPUT_BRAM_24_DMWIDTH/8-1:0] s_axis_bram_24_tstrb,
    input [C_INPUT_BRAM_24_DMWIDTH-1:0] s_axis_bram_24_tdata,
    output s_axis_bram_24_tready,
    input [C_INPUT_BRAM_24_ADDR_WIDTH-1:0] ap_bram_iarg_24_addr0,
    input [C_INPUT_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_din0,
    output [C_INPUT_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_dout0,
    input ap_bram_iarg_24_clk0,
    input ap_bram_iarg_24_rst0,
    input [C_INPUT_BRAM_24_WIDTH/8-1:0] ap_bram_iarg_24_we0,
    input ap_bram_iarg_24_en0,
    input [C_INPUT_BRAM_24_ADDR_WIDTH-1:0] ap_bram_iarg_24_addr1,
    input [C_INPUT_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_din1,
    output [C_INPUT_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_dout1,
    input ap_bram_iarg_24_clk1,
    input ap_bram_iarg_24_rst1,
    input [C_INPUT_BRAM_24_WIDTH/8-1:0] ap_bram_iarg_24_we1,
    input ap_bram_iarg_24_en1,
    //input AXI-Stream to BRAM interface 25
    input s_axis_bram_25_tlast,
    input s_axis_bram_25_tvalid,
    input [C_INPUT_BRAM_25_DMWIDTH/8-1:0] s_axis_bram_25_tkeep,
    input [C_INPUT_BRAM_25_DMWIDTH/8-1:0] s_axis_bram_25_tstrb,
    input [C_INPUT_BRAM_25_DMWIDTH-1:0] s_axis_bram_25_tdata,
    output s_axis_bram_25_tready,
    input [C_INPUT_BRAM_25_ADDR_WIDTH-1:0] ap_bram_iarg_25_addr0,
    input [C_INPUT_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_din0,
    output [C_INPUT_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_dout0,
    input ap_bram_iarg_25_clk0,
    input ap_bram_iarg_25_rst0,
    input [C_INPUT_BRAM_25_WIDTH/8-1:0] ap_bram_iarg_25_we0,
    input ap_bram_iarg_25_en0,
    input [C_INPUT_BRAM_25_ADDR_WIDTH-1:0] ap_bram_iarg_25_addr1,
    input [C_INPUT_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_din1,
    output [C_INPUT_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_dout1,
    input ap_bram_iarg_25_clk1,
    input ap_bram_iarg_25_rst1,
    input [C_INPUT_BRAM_25_WIDTH/8-1:0] ap_bram_iarg_25_we1,
    input ap_bram_iarg_25_en1,
    //input AXI-Stream to BRAM interface 26
    input s_axis_bram_26_tlast,
    input s_axis_bram_26_tvalid,
    input [C_INPUT_BRAM_26_DMWIDTH/8-1:0] s_axis_bram_26_tkeep,
    input [C_INPUT_BRAM_26_DMWIDTH/8-1:0] s_axis_bram_26_tstrb,
    input [C_INPUT_BRAM_26_DMWIDTH-1:0] s_axis_bram_26_tdata,
    output s_axis_bram_26_tready,
    input [C_INPUT_BRAM_26_ADDR_WIDTH-1:0] ap_bram_iarg_26_addr0,
    input [C_INPUT_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_din0,
    output [C_INPUT_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_dout0,
    input ap_bram_iarg_26_clk0,
    input ap_bram_iarg_26_rst0,
    input [C_INPUT_BRAM_26_WIDTH/8-1:0] ap_bram_iarg_26_we0,
    input ap_bram_iarg_26_en0,
    input [C_INPUT_BRAM_26_ADDR_WIDTH-1:0] ap_bram_iarg_26_addr1,
    input [C_INPUT_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_din1,
    output [C_INPUT_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_dout1,
    input ap_bram_iarg_26_clk1,
    input ap_bram_iarg_26_rst1,
    input [C_INPUT_BRAM_26_WIDTH/8-1:0] ap_bram_iarg_26_we1,
    input ap_bram_iarg_26_en1,
    //input AXI-Stream to BRAM interface 27
    input s_axis_bram_27_tlast,
    input s_axis_bram_27_tvalid,
    input [C_INPUT_BRAM_27_DMWIDTH/8-1:0] s_axis_bram_27_tkeep,
    input [C_INPUT_BRAM_27_DMWIDTH/8-1:0] s_axis_bram_27_tstrb,
    input [C_INPUT_BRAM_27_DMWIDTH-1:0] s_axis_bram_27_tdata,
    output s_axis_bram_27_tready,
    input [C_INPUT_BRAM_27_ADDR_WIDTH-1:0] ap_bram_iarg_27_addr0,
    input [C_INPUT_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_din0,
    output [C_INPUT_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_dout0,
    input ap_bram_iarg_27_clk0,
    input ap_bram_iarg_27_rst0,
    input [C_INPUT_BRAM_27_WIDTH/8-1:0] ap_bram_iarg_27_we0,
    input ap_bram_iarg_27_en0,
    input [C_INPUT_BRAM_27_ADDR_WIDTH-1:0] ap_bram_iarg_27_addr1,
    input [C_INPUT_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_din1,
    output [C_INPUT_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_dout1,
    input ap_bram_iarg_27_clk1,
    input ap_bram_iarg_27_rst1,
    input [C_INPUT_BRAM_27_WIDTH/8-1:0] ap_bram_iarg_27_we1,
    input ap_bram_iarg_27_en1,
    //input AXI-Stream to BRAM interface 28
    input s_axis_bram_28_tlast,
    input s_axis_bram_28_tvalid,
    input [C_INPUT_BRAM_28_DMWIDTH/8-1:0] s_axis_bram_28_tkeep,
    input [C_INPUT_BRAM_28_DMWIDTH/8-1:0] s_axis_bram_28_tstrb,
    input [C_INPUT_BRAM_28_DMWIDTH-1:0] s_axis_bram_28_tdata,
    output s_axis_bram_28_tready,
    input [C_INPUT_BRAM_28_ADDR_WIDTH-1:0] ap_bram_iarg_28_addr0,
    input [C_INPUT_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_din0,
    output [C_INPUT_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_dout0,
    input ap_bram_iarg_28_clk0,
    input ap_bram_iarg_28_rst0,
    input [C_INPUT_BRAM_28_WIDTH/8-1:0] ap_bram_iarg_28_we0,
    input ap_bram_iarg_28_en0,
    input [C_INPUT_BRAM_28_ADDR_WIDTH-1:0] ap_bram_iarg_28_addr1,
    input [C_INPUT_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_din1,
    output [C_INPUT_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_dout1,
    input ap_bram_iarg_28_clk1,
    input ap_bram_iarg_28_rst1,
    input [C_INPUT_BRAM_28_WIDTH/8-1:0] ap_bram_iarg_28_we1,
    input ap_bram_iarg_28_en1,
    //input AXI-Stream to BRAM interface 29
    input s_axis_bram_29_tlast,
    input s_axis_bram_29_tvalid,
    input [C_INPUT_BRAM_29_DMWIDTH/8-1:0] s_axis_bram_29_tkeep,
    input [C_INPUT_BRAM_29_DMWIDTH/8-1:0] s_axis_bram_29_tstrb,
    input [C_INPUT_BRAM_29_DMWIDTH-1:0] s_axis_bram_29_tdata,
    output s_axis_bram_29_tready,
    input [C_INPUT_BRAM_29_ADDR_WIDTH-1:0] ap_bram_iarg_29_addr0,
    input [C_INPUT_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_din0,
    output [C_INPUT_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_dout0,
    input ap_bram_iarg_29_clk0,
    input ap_bram_iarg_29_rst0,
    input [C_INPUT_BRAM_29_WIDTH/8-1:0] ap_bram_iarg_29_we0,
    input ap_bram_iarg_29_en0,
    input [C_INPUT_BRAM_29_ADDR_WIDTH-1:0] ap_bram_iarg_29_addr1,
    input [C_INPUT_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_din1,
    output [C_INPUT_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_dout1,
    input ap_bram_iarg_29_clk1,
    input ap_bram_iarg_29_rst1,
    input [C_INPUT_BRAM_29_WIDTH/8-1:0] ap_bram_iarg_29_we1,
    input ap_bram_iarg_29_en1,
    //input AXI-Stream to BRAM interface 30
    input s_axis_bram_30_tlast,
    input s_axis_bram_30_tvalid,
    input [C_INPUT_BRAM_30_DMWIDTH/8-1:0] s_axis_bram_30_tkeep,
    input [C_INPUT_BRAM_30_DMWIDTH/8-1:0] s_axis_bram_30_tstrb,
    input [C_INPUT_BRAM_30_DMWIDTH-1:0] s_axis_bram_30_tdata,
    output s_axis_bram_30_tready,
    input [C_INPUT_BRAM_30_ADDR_WIDTH-1:0] ap_bram_iarg_30_addr0,
    input [C_INPUT_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_din0,
    output [C_INPUT_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_dout0,
    input ap_bram_iarg_30_clk0,
    input ap_bram_iarg_30_rst0,
    input [C_INPUT_BRAM_30_WIDTH/8-1:0] ap_bram_iarg_30_we0,
    input ap_bram_iarg_30_en0,
    input [C_INPUT_BRAM_30_ADDR_WIDTH-1:0] ap_bram_iarg_30_addr1,
    input [C_INPUT_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_din1,
    output [C_INPUT_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_dout1,
    input ap_bram_iarg_30_clk1,
    input ap_bram_iarg_30_rst1,
    input [C_INPUT_BRAM_30_WIDTH/8-1:0] ap_bram_iarg_30_we1,
    input ap_bram_iarg_30_en1,
    //input AXI-Stream to BRAM interface 31
    input s_axis_bram_31_tlast,
    input s_axis_bram_31_tvalid,
    input [C_INPUT_BRAM_31_DMWIDTH/8-1:0] s_axis_bram_31_tkeep,
    input [C_INPUT_BRAM_31_DMWIDTH/8-1:0] s_axis_bram_31_tstrb,
    input [C_INPUT_BRAM_31_DMWIDTH-1:0] s_axis_bram_31_tdata,
    output s_axis_bram_31_tready,
    input [C_INPUT_BRAM_31_ADDR_WIDTH-1:0] ap_bram_iarg_31_addr0,
    input [C_INPUT_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_din0,
    output [C_INPUT_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_dout0,
    input ap_bram_iarg_31_clk0,
    input ap_bram_iarg_31_rst0,
    input [C_INPUT_BRAM_31_WIDTH/8-1:0] ap_bram_iarg_31_we0,
    input ap_bram_iarg_31_en0,
    input [C_INPUT_BRAM_31_ADDR_WIDTH-1:0] ap_bram_iarg_31_addr1,
    input [C_INPUT_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_din1,
    output [C_INPUT_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_dout1,
    input ap_bram_iarg_31_clk1,
    input ap_bram_iarg_31_rst1,
    input [C_INPUT_BRAM_31_WIDTH/8-1:0] ap_bram_iarg_31_we1,
    input ap_bram_iarg_31_en1,
    //input AXI-Stream to BRAM interface 32
    input s_axis_bram_32_tlast,
    input s_axis_bram_32_tvalid,
    input [C_INPUT_BRAM_32_DMWIDTH/8-1:0] s_axis_bram_32_tkeep,
    input [C_INPUT_BRAM_32_DMWIDTH/8-1:0] s_axis_bram_32_tstrb,
    input [C_INPUT_BRAM_32_DMWIDTH-1:0] s_axis_bram_32_tdata,
    output s_axis_bram_32_tready,
    input [C_INPUT_BRAM_32_ADDR_WIDTH-1:0] ap_bram_iarg_32_addr0,
    input [C_INPUT_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_din0,
    output [C_INPUT_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_dout0,
    input ap_bram_iarg_32_clk0,
    input ap_bram_iarg_32_rst0,
    input [C_INPUT_BRAM_32_WIDTH/8-1:0] ap_bram_iarg_32_we0,
    input ap_bram_iarg_32_en0,
    input [C_INPUT_BRAM_32_ADDR_WIDTH-1:0] ap_bram_iarg_32_addr1,
    input [C_INPUT_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_din1,
    output [C_INPUT_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_dout1,
    input ap_bram_iarg_32_clk1,
    input ap_bram_iarg_32_rst1,
    input [C_INPUT_BRAM_32_WIDTH/8-1:0] ap_bram_iarg_32_we1,
    input ap_bram_iarg_32_en1,
    //input AXI-Stream to BRAM interface 33
    input s_axis_bram_33_tlast,
    input s_axis_bram_33_tvalid,
    input [C_INPUT_BRAM_33_DMWIDTH/8-1:0] s_axis_bram_33_tkeep,
    input [C_INPUT_BRAM_33_DMWIDTH/8-1:0] s_axis_bram_33_tstrb,
    input [C_INPUT_BRAM_33_DMWIDTH-1:0] s_axis_bram_33_tdata,
    output s_axis_bram_33_tready,
    input [C_INPUT_BRAM_33_ADDR_WIDTH-1:0] ap_bram_iarg_33_addr0,
    input [C_INPUT_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_din0,
    output [C_INPUT_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_dout0,
    input ap_bram_iarg_33_clk0,
    input ap_bram_iarg_33_rst0,
    input [C_INPUT_BRAM_33_WIDTH/8-1:0] ap_bram_iarg_33_we0,
    input ap_bram_iarg_33_en0,
    input [C_INPUT_BRAM_33_ADDR_WIDTH-1:0] ap_bram_iarg_33_addr1,
    input [C_INPUT_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_din1,
    output [C_INPUT_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_dout1,
    input ap_bram_iarg_33_clk1,
    input ap_bram_iarg_33_rst1,
    input [C_INPUT_BRAM_33_WIDTH/8-1:0] ap_bram_iarg_33_we1,
    input ap_bram_iarg_33_en1,
    //input AXI-Stream to BRAM interface 34
    input s_axis_bram_34_tlast,
    input s_axis_bram_34_tvalid,
    input [C_INPUT_BRAM_34_DMWIDTH/8-1:0] s_axis_bram_34_tkeep,
    input [C_INPUT_BRAM_34_DMWIDTH/8-1:0] s_axis_bram_34_tstrb,
    input [C_INPUT_BRAM_34_DMWIDTH-1:0] s_axis_bram_34_tdata,
    output s_axis_bram_34_tready,
    input [C_INPUT_BRAM_34_ADDR_WIDTH-1:0] ap_bram_iarg_34_addr0,
    input [C_INPUT_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_din0,
    output [C_INPUT_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_dout0,
    input ap_bram_iarg_34_clk0,
    input ap_bram_iarg_34_rst0,
    input [C_INPUT_BRAM_34_WIDTH/8-1:0] ap_bram_iarg_34_we0,
    input ap_bram_iarg_34_en0,
    input [C_INPUT_BRAM_34_ADDR_WIDTH-1:0] ap_bram_iarg_34_addr1,
    input [C_INPUT_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_din1,
    output [C_INPUT_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_dout1,
    input ap_bram_iarg_34_clk1,
    input ap_bram_iarg_34_rst1,
    input [C_INPUT_BRAM_34_WIDTH/8-1:0] ap_bram_iarg_34_we1,
    input ap_bram_iarg_34_en1,
    //input AXI-Stream to BRAM interface 35
    input s_axis_bram_35_tlast,
    input s_axis_bram_35_tvalid,
    input [C_INPUT_BRAM_35_DMWIDTH/8-1:0] s_axis_bram_35_tkeep,
    input [C_INPUT_BRAM_35_DMWIDTH/8-1:0] s_axis_bram_35_tstrb,
    input [C_INPUT_BRAM_35_DMWIDTH-1:0] s_axis_bram_35_tdata,
    output s_axis_bram_35_tready,
    input [C_INPUT_BRAM_35_ADDR_WIDTH-1:0] ap_bram_iarg_35_addr0,
    input [C_INPUT_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_din0,
    output [C_INPUT_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_dout0,
    input ap_bram_iarg_35_clk0,
    input ap_bram_iarg_35_rst0,
    input [C_INPUT_BRAM_35_WIDTH/8-1:0] ap_bram_iarg_35_we0,
    input ap_bram_iarg_35_en0,
    input [C_INPUT_BRAM_35_ADDR_WIDTH-1:0] ap_bram_iarg_35_addr1,
    input [C_INPUT_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_din1,
    output [C_INPUT_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_dout1,
    input ap_bram_iarg_35_clk1,
    input ap_bram_iarg_35_rst1,
    input [C_INPUT_BRAM_35_WIDTH/8-1:0] ap_bram_iarg_35_we1,
    input ap_bram_iarg_35_en1,
    //input AXI-Stream to BRAM interface 36
    input s_axis_bram_36_tlast,
    input s_axis_bram_36_tvalid,
    input [C_INPUT_BRAM_36_DMWIDTH/8-1:0] s_axis_bram_36_tkeep,
    input [C_INPUT_BRAM_36_DMWIDTH/8-1:0] s_axis_bram_36_tstrb,
    input [C_INPUT_BRAM_36_DMWIDTH-1:0] s_axis_bram_36_tdata,
    output s_axis_bram_36_tready,
    input [C_INPUT_BRAM_36_ADDR_WIDTH-1:0] ap_bram_iarg_36_addr0,
    input [C_INPUT_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_din0,
    output [C_INPUT_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_dout0,
    input ap_bram_iarg_36_clk0,
    input ap_bram_iarg_36_rst0,
    input [C_INPUT_BRAM_36_WIDTH/8-1:0] ap_bram_iarg_36_we0,
    input ap_bram_iarg_36_en0,
    input [C_INPUT_BRAM_36_ADDR_WIDTH-1:0] ap_bram_iarg_36_addr1,
    input [C_INPUT_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_din1,
    output [C_INPUT_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_dout1,
    input ap_bram_iarg_36_clk1,
    input ap_bram_iarg_36_rst1,
    input [C_INPUT_BRAM_36_WIDTH/8-1:0] ap_bram_iarg_36_we1,
    input ap_bram_iarg_36_en1,
    //input AXI-Stream to BRAM interface 37
    input s_axis_bram_37_tlast,
    input s_axis_bram_37_tvalid,
    input [C_INPUT_BRAM_37_DMWIDTH/8-1:0] s_axis_bram_37_tkeep,
    input [C_INPUT_BRAM_37_DMWIDTH/8-1:0] s_axis_bram_37_tstrb,
    input [C_INPUT_BRAM_37_DMWIDTH-1:0] s_axis_bram_37_tdata,
    output s_axis_bram_37_tready,
    input [C_INPUT_BRAM_37_ADDR_WIDTH-1:0] ap_bram_iarg_37_addr0,
    input [C_INPUT_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_din0,
    output [C_INPUT_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_dout0,
    input ap_bram_iarg_37_clk0,
    input ap_bram_iarg_37_rst0,
    input [C_INPUT_BRAM_37_WIDTH/8-1:0] ap_bram_iarg_37_we0,
    input ap_bram_iarg_37_en0,
    input [C_INPUT_BRAM_37_ADDR_WIDTH-1:0] ap_bram_iarg_37_addr1,
    input [C_INPUT_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_din1,
    output [C_INPUT_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_dout1,
    input ap_bram_iarg_37_clk1,
    input ap_bram_iarg_37_rst1,
    input [C_INPUT_BRAM_37_WIDTH/8-1:0] ap_bram_iarg_37_we1,
    input ap_bram_iarg_37_en1,
    //input AXI-Stream to BRAM interface 38
    input s_axis_bram_38_tlast,
    input s_axis_bram_38_tvalid,
    input [C_INPUT_BRAM_38_DMWIDTH/8-1:0] s_axis_bram_38_tkeep,
    input [C_INPUT_BRAM_38_DMWIDTH/8-1:0] s_axis_bram_38_tstrb,
    input [C_INPUT_BRAM_38_DMWIDTH-1:0] s_axis_bram_38_tdata,
    output s_axis_bram_38_tready,
    input [C_INPUT_BRAM_38_ADDR_WIDTH-1:0] ap_bram_iarg_38_addr0,
    input [C_INPUT_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_din0,
    output [C_INPUT_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_dout0,
    input ap_bram_iarg_38_clk0,
    input ap_bram_iarg_38_rst0,
    input [C_INPUT_BRAM_38_WIDTH/8-1:0] ap_bram_iarg_38_we0,
    input ap_bram_iarg_38_en0,
    input [C_INPUT_BRAM_38_ADDR_WIDTH-1:0] ap_bram_iarg_38_addr1,
    input [C_INPUT_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_din1,
    output [C_INPUT_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_dout1,
    input ap_bram_iarg_38_clk1,
    input ap_bram_iarg_38_rst1,
    input [C_INPUT_BRAM_38_WIDTH/8-1:0] ap_bram_iarg_38_we1,
    input ap_bram_iarg_38_en1,
    //input AXI-Stream to BRAM interface 39
    input s_axis_bram_39_tlast,
    input s_axis_bram_39_tvalid,
    input [C_INPUT_BRAM_39_DMWIDTH/8-1:0] s_axis_bram_39_tkeep,
    input [C_INPUT_BRAM_39_DMWIDTH/8-1:0] s_axis_bram_39_tstrb,
    input [C_INPUT_BRAM_39_DMWIDTH-1:0] s_axis_bram_39_tdata,
    output s_axis_bram_39_tready,
    input [C_INPUT_BRAM_39_ADDR_WIDTH-1:0] ap_bram_iarg_39_addr0,
    input [C_INPUT_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_din0,
    output [C_INPUT_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_dout0,
    input ap_bram_iarg_39_clk0,
    input ap_bram_iarg_39_rst0,
    input [C_INPUT_BRAM_39_WIDTH/8-1:0] ap_bram_iarg_39_we0,
    input ap_bram_iarg_39_en0,
    input [C_INPUT_BRAM_39_ADDR_WIDTH-1:0] ap_bram_iarg_39_addr1,
    input [C_INPUT_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_din1,
    output [C_INPUT_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_dout1,
    input ap_bram_iarg_39_clk1,
    input ap_bram_iarg_39_rst1,
    input [C_INPUT_BRAM_39_WIDTH/8-1:0] ap_bram_iarg_39_we1,
    input ap_bram_iarg_39_en1,
    //input AXI-Stream to BRAM interface 40
    input s_axis_bram_40_tlast,
    input s_axis_bram_40_tvalid,
    input [C_INPUT_BRAM_40_DMWIDTH/8-1:0] s_axis_bram_40_tkeep,
    input [C_INPUT_BRAM_40_DMWIDTH/8-1:0] s_axis_bram_40_tstrb,
    input [C_INPUT_BRAM_40_DMWIDTH-1:0] s_axis_bram_40_tdata,
    output s_axis_bram_40_tready,
    input [C_INPUT_BRAM_40_ADDR_WIDTH-1:0] ap_bram_iarg_40_addr0,
    input [C_INPUT_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_din0,
    output [C_INPUT_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_dout0,
    input ap_bram_iarg_40_clk0,
    input ap_bram_iarg_40_rst0,
    input [C_INPUT_BRAM_40_WIDTH/8-1:0] ap_bram_iarg_40_we0,
    input ap_bram_iarg_40_en0,
    input [C_INPUT_BRAM_40_ADDR_WIDTH-1:0] ap_bram_iarg_40_addr1,
    input [C_INPUT_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_din1,
    output [C_INPUT_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_dout1,
    input ap_bram_iarg_40_clk1,
    input ap_bram_iarg_40_rst1,
    input [C_INPUT_BRAM_40_WIDTH/8-1:0] ap_bram_iarg_40_we1,
    input ap_bram_iarg_40_en1,
    //input AXI-Stream to BRAM interface 41
    input s_axis_bram_41_tlast,
    input s_axis_bram_41_tvalid,
    input [C_INPUT_BRAM_41_DMWIDTH/8-1:0] s_axis_bram_41_tkeep,
    input [C_INPUT_BRAM_41_DMWIDTH/8-1:0] s_axis_bram_41_tstrb,
    input [C_INPUT_BRAM_41_DMWIDTH-1:0] s_axis_bram_41_tdata,
    output s_axis_bram_41_tready,
    input [C_INPUT_BRAM_41_ADDR_WIDTH-1:0] ap_bram_iarg_41_addr0,
    input [C_INPUT_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_din0,
    output [C_INPUT_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_dout0,
    input ap_bram_iarg_41_clk0,
    input ap_bram_iarg_41_rst0,
    input [C_INPUT_BRAM_41_WIDTH/8-1:0] ap_bram_iarg_41_we0,
    input ap_bram_iarg_41_en0,
    input [C_INPUT_BRAM_41_ADDR_WIDTH-1:0] ap_bram_iarg_41_addr1,
    input [C_INPUT_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_din1,
    output [C_INPUT_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_dout1,
    input ap_bram_iarg_41_clk1,
    input ap_bram_iarg_41_rst1,
    input [C_INPUT_BRAM_41_WIDTH/8-1:0] ap_bram_iarg_41_we1,
    input ap_bram_iarg_41_en1,
    //input AXI-Stream to BRAM interface 42
    input s_axis_bram_42_tlast,
    input s_axis_bram_42_tvalid,
    input [C_INPUT_BRAM_42_DMWIDTH/8-1:0] s_axis_bram_42_tkeep,
    input [C_INPUT_BRAM_42_DMWIDTH/8-1:0] s_axis_bram_42_tstrb,
    input [C_INPUT_BRAM_42_DMWIDTH-1:0] s_axis_bram_42_tdata,
    output s_axis_bram_42_tready,
    input [C_INPUT_BRAM_42_ADDR_WIDTH-1:0] ap_bram_iarg_42_addr0,
    input [C_INPUT_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_din0,
    output [C_INPUT_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_dout0,
    input ap_bram_iarg_42_clk0,
    input ap_bram_iarg_42_rst0,
    input [C_INPUT_BRAM_42_WIDTH/8-1:0] ap_bram_iarg_42_we0,
    input ap_bram_iarg_42_en0,
    input [C_INPUT_BRAM_42_ADDR_WIDTH-1:0] ap_bram_iarg_42_addr1,
    input [C_INPUT_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_din1,
    output [C_INPUT_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_dout1,
    input ap_bram_iarg_42_clk1,
    input ap_bram_iarg_42_rst1,
    input [C_INPUT_BRAM_42_WIDTH/8-1:0] ap_bram_iarg_42_we1,
    input ap_bram_iarg_42_en1,
    //input AXI-Stream to BRAM interface 43
    input s_axis_bram_43_tlast,
    input s_axis_bram_43_tvalid,
    input [C_INPUT_BRAM_43_DMWIDTH/8-1:0] s_axis_bram_43_tkeep,
    input [C_INPUT_BRAM_43_DMWIDTH/8-1:0] s_axis_bram_43_tstrb,
    input [C_INPUT_BRAM_43_DMWIDTH-1:0] s_axis_bram_43_tdata,
    output s_axis_bram_43_tready,
    input [C_INPUT_BRAM_43_ADDR_WIDTH-1:0] ap_bram_iarg_43_addr0,
    input [C_INPUT_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_din0,
    output [C_INPUT_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_dout0,
    input ap_bram_iarg_43_clk0,
    input ap_bram_iarg_43_rst0,
    input [C_INPUT_BRAM_43_WIDTH/8-1:0] ap_bram_iarg_43_we0,
    input ap_bram_iarg_43_en0,
    input [C_INPUT_BRAM_43_ADDR_WIDTH-1:0] ap_bram_iarg_43_addr1,
    input [C_INPUT_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_din1,
    output [C_INPUT_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_dout1,
    input ap_bram_iarg_43_clk1,
    input ap_bram_iarg_43_rst1,
    input [C_INPUT_BRAM_43_WIDTH/8-1:0] ap_bram_iarg_43_we1,
    input ap_bram_iarg_43_en1,
    //input AXI-Stream to BRAM interface 44
    input s_axis_bram_44_tlast,
    input s_axis_bram_44_tvalid,
    input [C_INPUT_BRAM_44_DMWIDTH/8-1:0] s_axis_bram_44_tkeep,
    input [C_INPUT_BRAM_44_DMWIDTH/8-1:0] s_axis_bram_44_tstrb,
    input [C_INPUT_BRAM_44_DMWIDTH-1:0] s_axis_bram_44_tdata,
    output s_axis_bram_44_tready,
    input [C_INPUT_BRAM_44_ADDR_WIDTH-1:0] ap_bram_iarg_44_addr0,
    input [C_INPUT_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_din0,
    output [C_INPUT_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_dout0,
    input ap_bram_iarg_44_clk0,
    input ap_bram_iarg_44_rst0,
    input [C_INPUT_BRAM_44_WIDTH/8-1:0] ap_bram_iarg_44_we0,
    input ap_bram_iarg_44_en0,
    input [C_INPUT_BRAM_44_ADDR_WIDTH-1:0] ap_bram_iarg_44_addr1,
    input [C_INPUT_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_din1,
    output [C_INPUT_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_dout1,
    input ap_bram_iarg_44_clk1,
    input ap_bram_iarg_44_rst1,
    input [C_INPUT_BRAM_44_WIDTH/8-1:0] ap_bram_iarg_44_we1,
    input ap_bram_iarg_44_en1,
    //input AXI-Stream to BRAM interface 45
    input s_axis_bram_45_tlast,
    input s_axis_bram_45_tvalid,
    input [C_INPUT_BRAM_45_DMWIDTH/8-1:0] s_axis_bram_45_tkeep,
    input [C_INPUT_BRAM_45_DMWIDTH/8-1:0] s_axis_bram_45_tstrb,
    input [C_INPUT_BRAM_45_DMWIDTH-1:0] s_axis_bram_45_tdata,
    output s_axis_bram_45_tready,
    input [C_INPUT_BRAM_45_ADDR_WIDTH-1:0] ap_bram_iarg_45_addr0,
    input [C_INPUT_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_din0,
    output [C_INPUT_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_dout0,
    input ap_bram_iarg_45_clk0,
    input ap_bram_iarg_45_rst0,
    input [C_INPUT_BRAM_45_WIDTH/8-1:0] ap_bram_iarg_45_we0,
    input ap_bram_iarg_45_en0,
    input [C_INPUT_BRAM_45_ADDR_WIDTH-1:0] ap_bram_iarg_45_addr1,
    input [C_INPUT_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_din1,
    output [C_INPUT_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_dout1,
    input ap_bram_iarg_45_clk1,
    input ap_bram_iarg_45_rst1,
    input [C_INPUT_BRAM_45_WIDTH/8-1:0] ap_bram_iarg_45_we1,
    input ap_bram_iarg_45_en1,
    //input AXI-Stream to BRAM interface 46
    input s_axis_bram_46_tlast,
    input s_axis_bram_46_tvalid,
    input [C_INPUT_BRAM_46_DMWIDTH/8-1:0] s_axis_bram_46_tkeep,
    input [C_INPUT_BRAM_46_DMWIDTH/8-1:0] s_axis_bram_46_tstrb,
    input [C_INPUT_BRAM_46_DMWIDTH-1:0] s_axis_bram_46_tdata,
    output s_axis_bram_46_tready,
    input [C_INPUT_BRAM_46_ADDR_WIDTH-1:0] ap_bram_iarg_46_addr0,
    input [C_INPUT_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_din0,
    output [C_INPUT_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_dout0,
    input ap_bram_iarg_46_clk0,
    input ap_bram_iarg_46_rst0,
    input [C_INPUT_BRAM_46_WIDTH/8-1:0] ap_bram_iarg_46_we0,
    input ap_bram_iarg_46_en0,
    input [C_INPUT_BRAM_46_ADDR_WIDTH-1:0] ap_bram_iarg_46_addr1,
    input [C_INPUT_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_din1,
    output [C_INPUT_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_dout1,
    input ap_bram_iarg_46_clk1,
    input ap_bram_iarg_46_rst1,
    input [C_INPUT_BRAM_46_WIDTH/8-1:0] ap_bram_iarg_46_we1,
    input ap_bram_iarg_46_en1,
    //input AXI-Stream to BRAM interface 47
    input s_axis_bram_47_tlast,
    input s_axis_bram_47_tvalid,
    input [C_INPUT_BRAM_47_DMWIDTH/8-1:0] s_axis_bram_47_tkeep,
    input [C_INPUT_BRAM_47_DMWIDTH/8-1:0] s_axis_bram_47_tstrb,
    input [C_INPUT_BRAM_47_DMWIDTH-1:0] s_axis_bram_47_tdata,
    output s_axis_bram_47_tready,
    input [C_INPUT_BRAM_47_ADDR_WIDTH-1:0] ap_bram_iarg_47_addr0,
    input [C_INPUT_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_din0,
    output [C_INPUT_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_dout0,
    input ap_bram_iarg_47_clk0,
    input ap_bram_iarg_47_rst0,
    input [C_INPUT_BRAM_47_WIDTH/8-1:0] ap_bram_iarg_47_we0,
    input ap_bram_iarg_47_en0,
    input [C_INPUT_BRAM_47_ADDR_WIDTH-1:0] ap_bram_iarg_47_addr1,
    input [C_INPUT_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_din1,
    output [C_INPUT_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_dout1,
    input ap_bram_iarg_47_clk1,
    input ap_bram_iarg_47_rst1,
    input [C_INPUT_BRAM_47_WIDTH/8-1:0] ap_bram_iarg_47_we1,
    input ap_bram_iarg_47_en1,
    //input AXI-Stream to BRAM interface 48
    input s_axis_bram_48_tlast,
    input s_axis_bram_48_tvalid,
    input [C_INPUT_BRAM_48_DMWIDTH/8-1:0] s_axis_bram_48_tkeep,
    input [C_INPUT_BRAM_48_DMWIDTH/8-1:0] s_axis_bram_48_tstrb,
    input [C_INPUT_BRAM_48_DMWIDTH-1:0] s_axis_bram_48_tdata,
    output s_axis_bram_48_tready,
    input [C_INPUT_BRAM_48_ADDR_WIDTH-1:0] ap_bram_iarg_48_addr0,
    input [C_INPUT_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_din0,
    output [C_INPUT_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_dout0,
    input ap_bram_iarg_48_clk0,
    input ap_bram_iarg_48_rst0,
    input [C_INPUT_BRAM_48_WIDTH/8-1:0] ap_bram_iarg_48_we0,
    input ap_bram_iarg_48_en0,
    input [C_INPUT_BRAM_48_ADDR_WIDTH-1:0] ap_bram_iarg_48_addr1,
    input [C_INPUT_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_din1,
    output [C_INPUT_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_dout1,
    input ap_bram_iarg_48_clk1,
    input ap_bram_iarg_48_rst1,
    input [C_INPUT_BRAM_48_WIDTH/8-1:0] ap_bram_iarg_48_we1,
    input ap_bram_iarg_48_en1,
    //input AXI-Stream to BRAM interface 49
    input s_axis_bram_49_tlast,
    input s_axis_bram_49_tvalid,
    input [C_INPUT_BRAM_49_DMWIDTH/8-1:0] s_axis_bram_49_tkeep,
    input [C_INPUT_BRAM_49_DMWIDTH/8-1:0] s_axis_bram_49_tstrb,
    input [C_INPUT_BRAM_49_DMWIDTH-1:0] s_axis_bram_49_tdata,
    output s_axis_bram_49_tready,
    input [C_INPUT_BRAM_49_ADDR_WIDTH-1:0] ap_bram_iarg_49_addr0,
    input [C_INPUT_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_din0,
    output [C_INPUT_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_dout0,
    input ap_bram_iarg_49_clk0,
    input ap_bram_iarg_49_rst0,
    input [C_INPUT_BRAM_49_WIDTH/8-1:0] ap_bram_iarg_49_we0,
    input ap_bram_iarg_49_en0,
    input [C_INPUT_BRAM_49_ADDR_WIDTH-1:0] ap_bram_iarg_49_addr1,
    input [C_INPUT_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_din1,
    output [C_INPUT_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_dout1,
    input ap_bram_iarg_49_clk1,
    input ap_bram_iarg_49_rst1,
    input [C_INPUT_BRAM_49_WIDTH/8-1:0] ap_bram_iarg_49_we1,
    input ap_bram_iarg_49_en1,
    //input AXI-Stream to BRAM interface 50
    input s_axis_bram_50_tlast,
    input s_axis_bram_50_tvalid,
    input [C_INPUT_BRAM_50_DMWIDTH/8-1:0] s_axis_bram_50_tkeep,
    input [C_INPUT_BRAM_50_DMWIDTH/8-1:0] s_axis_bram_50_tstrb,
    input [C_INPUT_BRAM_50_DMWIDTH-1:0] s_axis_bram_50_tdata,
    output s_axis_bram_50_tready,
    input [C_INPUT_BRAM_50_ADDR_WIDTH-1:0] ap_bram_iarg_50_addr0,
    input [C_INPUT_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_din0,
    output [C_INPUT_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_dout0,
    input ap_bram_iarg_50_clk0,
    input ap_bram_iarg_50_rst0,
    input [C_INPUT_BRAM_50_WIDTH/8-1:0] ap_bram_iarg_50_we0,
    input ap_bram_iarg_50_en0,
    input [C_INPUT_BRAM_50_ADDR_WIDTH-1:0] ap_bram_iarg_50_addr1,
    input [C_INPUT_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_din1,
    output [C_INPUT_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_dout1,
    input ap_bram_iarg_50_clk1,
    input ap_bram_iarg_50_rst1,
    input [C_INPUT_BRAM_50_WIDTH/8-1:0] ap_bram_iarg_50_we1,
    input ap_bram_iarg_50_en1,
    //input AXI-Stream to BRAM interface 51
    input s_axis_bram_51_tlast,
    input s_axis_bram_51_tvalid,
    input [C_INPUT_BRAM_51_DMWIDTH/8-1:0] s_axis_bram_51_tkeep,
    input [C_INPUT_BRAM_51_DMWIDTH/8-1:0] s_axis_bram_51_tstrb,
    input [C_INPUT_BRAM_51_DMWIDTH-1:0] s_axis_bram_51_tdata,
    output s_axis_bram_51_tready,
    input [C_INPUT_BRAM_51_ADDR_WIDTH-1:0] ap_bram_iarg_51_addr0,
    input [C_INPUT_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_din0,
    output [C_INPUT_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_dout0,
    input ap_bram_iarg_51_clk0,
    input ap_bram_iarg_51_rst0,
    input [C_INPUT_BRAM_51_WIDTH/8-1:0] ap_bram_iarg_51_we0,
    input ap_bram_iarg_51_en0,
    input [C_INPUT_BRAM_51_ADDR_WIDTH-1:0] ap_bram_iarg_51_addr1,
    input [C_INPUT_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_din1,
    output [C_INPUT_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_dout1,
    input ap_bram_iarg_51_clk1,
    input ap_bram_iarg_51_rst1,
    input [C_INPUT_BRAM_51_WIDTH/8-1:0] ap_bram_iarg_51_we1,
    input ap_bram_iarg_51_en1,
    //input AXI-Stream to BRAM interface 52
    input s_axis_bram_52_tlast,
    input s_axis_bram_52_tvalid,
    input [C_INPUT_BRAM_52_DMWIDTH/8-1:0] s_axis_bram_52_tkeep,
    input [C_INPUT_BRAM_52_DMWIDTH/8-1:0] s_axis_bram_52_tstrb,
    input [C_INPUT_BRAM_52_DMWIDTH-1:0] s_axis_bram_52_tdata,
    output s_axis_bram_52_tready,
    input [C_INPUT_BRAM_52_ADDR_WIDTH-1:0] ap_bram_iarg_52_addr0,
    input [C_INPUT_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_din0,
    output [C_INPUT_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_dout0,
    input ap_bram_iarg_52_clk0,
    input ap_bram_iarg_52_rst0,
    input [C_INPUT_BRAM_52_WIDTH/8-1:0] ap_bram_iarg_52_we0,
    input ap_bram_iarg_52_en0,
    input [C_INPUT_BRAM_52_ADDR_WIDTH-1:0] ap_bram_iarg_52_addr1,
    input [C_INPUT_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_din1,
    output [C_INPUT_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_dout1,
    input ap_bram_iarg_52_clk1,
    input ap_bram_iarg_52_rst1,
    input [C_INPUT_BRAM_52_WIDTH/8-1:0] ap_bram_iarg_52_we1,
    input ap_bram_iarg_52_en1,
    //input AXI-Stream to BRAM interface 53
    input s_axis_bram_53_tlast,
    input s_axis_bram_53_tvalid,
    input [C_INPUT_BRAM_53_DMWIDTH/8-1:0] s_axis_bram_53_tkeep,
    input [C_INPUT_BRAM_53_DMWIDTH/8-1:0] s_axis_bram_53_tstrb,
    input [C_INPUT_BRAM_53_DMWIDTH-1:0] s_axis_bram_53_tdata,
    output s_axis_bram_53_tready,
    input [C_INPUT_BRAM_53_ADDR_WIDTH-1:0] ap_bram_iarg_53_addr0,
    input [C_INPUT_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_din0,
    output [C_INPUT_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_dout0,
    input ap_bram_iarg_53_clk0,
    input ap_bram_iarg_53_rst0,
    input [C_INPUT_BRAM_53_WIDTH/8-1:0] ap_bram_iarg_53_we0,
    input ap_bram_iarg_53_en0,
    input [C_INPUT_BRAM_53_ADDR_WIDTH-1:0] ap_bram_iarg_53_addr1,
    input [C_INPUT_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_din1,
    output [C_INPUT_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_dout1,
    input ap_bram_iarg_53_clk1,
    input ap_bram_iarg_53_rst1,
    input [C_INPUT_BRAM_53_WIDTH/8-1:0] ap_bram_iarg_53_we1,
    input ap_bram_iarg_53_en1,
    //input AXI-Stream to BRAM interface 54
    input s_axis_bram_54_tlast,
    input s_axis_bram_54_tvalid,
    input [C_INPUT_BRAM_54_DMWIDTH/8-1:0] s_axis_bram_54_tkeep,
    input [C_INPUT_BRAM_54_DMWIDTH/8-1:0] s_axis_bram_54_tstrb,
    input [C_INPUT_BRAM_54_DMWIDTH-1:0] s_axis_bram_54_tdata,
    output s_axis_bram_54_tready,
    input [C_INPUT_BRAM_54_ADDR_WIDTH-1:0] ap_bram_iarg_54_addr0,
    input [C_INPUT_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_din0,
    output [C_INPUT_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_dout0,
    input ap_bram_iarg_54_clk0,
    input ap_bram_iarg_54_rst0,
    input [C_INPUT_BRAM_54_WIDTH/8-1:0] ap_bram_iarg_54_we0,
    input ap_bram_iarg_54_en0,
    input [C_INPUT_BRAM_54_ADDR_WIDTH-1:0] ap_bram_iarg_54_addr1,
    input [C_INPUT_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_din1,
    output [C_INPUT_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_dout1,
    input ap_bram_iarg_54_clk1,
    input ap_bram_iarg_54_rst1,
    input [C_INPUT_BRAM_54_WIDTH/8-1:0] ap_bram_iarg_54_we1,
    input ap_bram_iarg_54_en1,
    //input AXI-Stream to BRAM interface 55
    input s_axis_bram_55_tlast,
    input s_axis_bram_55_tvalid,
    input [C_INPUT_BRAM_55_DMWIDTH/8-1:0] s_axis_bram_55_tkeep,
    input [C_INPUT_BRAM_55_DMWIDTH/8-1:0] s_axis_bram_55_tstrb,
    input [C_INPUT_BRAM_55_DMWIDTH-1:0] s_axis_bram_55_tdata,
    output s_axis_bram_55_tready,
    input [C_INPUT_BRAM_55_ADDR_WIDTH-1:0] ap_bram_iarg_55_addr0,
    input [C_INPUT_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_din0,
    output [C_INPUT_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_dout0,
    input ap_bram_iarg_55_clk0,
    input ap_bram_iarg_55_rst0,
    input [C_INPUT_BRAM_55_WIDTH/8-1:0] ap_bram_iarg_55_we0,
    input ap_bram_iarg_55_en0,
    input [C_INPUT_BRAM_55_ADDR_WIDTH-1:0] ap_bram_iarg_55_addr1,
    input [C_INPUT_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_din1,
    output [C_INPUT_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_dout1,
    input ap_bram_iarg_55_clk1,
    input ap_bram_iarg_55_rst1,
    input [C_INPUT_BRAM_55_WIDTH/8-1:0] ap_bram_iarg_55_we1,
    input ap_bram_iarg_55_en1,
    //input AXI-Stream to BRAM interface 56
    input s_axis_bram_56_tlast,
    input s_axis_bram_56_tvalid,
    input [C_INPUT_BRAM_56_DMWIDTH/8-1:0] s_axis_bram_56_tkeep,
    input [C_INPUT_BRAM_56_DMWIDTH/8-1:0] s_axis_bram_56_tstrb,
    input [C_INPUT_BRAM_56_DMWIDTH-1:0] s_axis_bram_56_tdata,
    output s_axis_bram_56_tready,
    input [C_INPUT_BRAM_56_ADDR_WIDTH-1:0] ap_bram_iarg_56_addr0,
    input [C_INPUT_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_din0,
    output [C_INPUT_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_dout0,
    input ap_bram_iarg_56_clk0,
    input ap_bram_iarg_56_rst0,
    input [C_INPUT_BRAM_56_WIDTH/8-1:0] ap_bram_iarg_56_we0,
    input ap_bram_iarg_56_en0,
    input [C_INPUT_BRAM_56_ADDR_WIDTH-1:0] ap_bram_iarg_56_addr1,
    input [C_INPUT_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_din1,
    output [C_INPUT_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_dout1,
    input ap_bram_iarg_56_clk1,
    input ap_bram_iarg_56_rst1,
    input [C_INPUT_BRAM_56_WIDTH/8-1:0] ap_bram_iarg_56_we1,
    input ap_bram_iarg_56_en1,
    //input AXI-Stream to BRAM interface 57
    input s_axis_bram_57_tlast,
    input s_axis_bram_57_tvalid,
    input [C_INPUT_BRAM_57_DMWIDTH/8-1:0] s_axis_bram_57_tkeep,
    input [C_INPUT_BRAM_57_DMWIDTH/8-1:0] s_axis_bram_57_tstrb,
    input [C_INPUT_BRAM_57_DMWIDTH-1:0] s_axis_bram_57_tdata,
    output s_axis_bram_57_tready,
    input [C_INPUT_BRAM_57_ADDR_WIDTH-1:0] ap_bram_iarg_57_addr0,
    input [C_INPUT_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_din0,
    output [C_INPUT_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_dout0,
    input ap_bram_iarg_57_clk0,
    input ap_bram_iarg_57_rst0,
    input [C_INPUT_BRAM_57_WIDTH/8-1:0] ap_bram_iarg_57_we0,
    input ap_bram_iarg_57_en0,
    input [C_INPUT_BRAM_57_ADDR_WIDTH-1:0] ap_bram_iarg_57_addr1,
    input [C_INPUT_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_din1,
    output [C_INPUT_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_dout1,
    input ap_bram_iarg_57_clk1,
    input ap_bram_iarg_57_rst1,
    input [C_INPUT_BRAM_57_WIDTH/8-1:0] ap_bram_iarg_57_we1,
    input ap_bram_iarg_57_en1,
    //input AXI-Stream to BRAM interface 58
    input s_axis_bram_58_tlast,
    input s_axis_bram_58_tvalid,
    input [C_INPUT_BRAM_58_DMWIDTH/8-1:0] s_axis_bram_58_tkeep,
    input [C_INPUT_BRAM_58_DMWIDTH/8-1:0] s_axis_bram_58_tstrb,
    input [C_INPUT_BRAM_58_DMWIDTH-1:0] s_axis_bram_58_tdata,
    output s_axis_bram_58_tready,
    input [C_INPUT_BRAM_58_ADDR_WIDTH-1:0] ap_bram_iarg_58_addr0,
    input [C_INPUT_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_din0,
    output [C_INPUT_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_dout0,
    input ap_bram_iarg_58_clk0,
    input ap_bram_iarg_58_rst0,
    input [C_INPUT_BRAM_58_WIDTH/8-1:0] ap_bram_iarg_58_we0,
    input ap_bram_iarg_58_en0,
    input [C_INPUT_BRAM_58_ADDR_WIDTH-1:0] ap_bram_iarg_58_addr1,
    input [C_INPUT_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_din1,
    output [C_INPUT_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_dout1,
    input ap_bram_iarg_58_clk1,
    input ap_bram_iarg_58_rst1,
    input [C_INPUT_BRAM_58_WIDTH/8-1:0] ap_bram_iarg_58_we1,
    input ap_bram_iarg_58_en1,
    //input AXI-Stream to BRAM interface 59
    input s_axis_bram_59_tlast,
    input s_axis_bram_59_tvalid,
    input [C_INPUT_BRAM_59_DMWIDTH/8-1:0] s_axis_bram_59_tkeep,
    input [C_INPUT_BRAM_59_DMWIDTH/8-1:0] s_axis_bram_59_tstrb,
    input [C_INPUT_BRAM_59_DMWIDTH-1:0] s_axis_bram_59_tdata,
    output s_axis_bram_59_tready,
    input [C_INPUT_BRAM_59_ADDR_WIDTH-1:0] ap_bram_iarg_59_addr0,
    input [C_INPUT_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_din0,
    output [C_INPUT_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_dout0,
    input ap_bram_iarg_59_clk0,
    input ap_bram_iarg_59_rst0,
    input [C_INPUT_BRAM_59_WIDTH/8-1:0] ap_bram_iarg_59_we0,
    input ap_bram_iarg_59_en0,
    input [C_INPUT_BRAM_59_ADDR_WIDTH-1:0] ap_bram_iarg_59_addr1,
    input [C_INPUT_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_din1,
    output [C_INPUT_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_dout1,
    input ap_bram_iarg_59_clk1,
    input ap_bram_iarg_59_rst1,
    input [C_INPUT_BRAM_59_WIDTH/8-1:0] ap_bram_iarg_59_we1,
    input ap_bram_iarg_59_en1,
    //input AXI-Stream to BRAM interface 60
    input s_axis_bram_60_tlast,
    input s_axis_bram_60_tvalid,
    input [C_INPUT_BRAM_60_DMWIDTH/8-1:0] s_axis_bram_60_tkeep,
    input [C_INPUT_BRAM_60_DMWIDTH/8-1:0] s_axis_bram_60_tstrb,
    input [C_INPUT_BRAM_60_DMWIDTH-1:0] s_axis_bram_60_tdata,
    output s_axis_bram_60_tready,
    input [C_INPUT_BRAM_60_ADDR_WIDTH-1:0] ap_bram_iarg_60_addr0,
    input [C_INPUT_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_din0,
    output [C_INPUT_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_dout0,
    input ap_bram_iarg_60_clk0,
    input ap_bram_iarg_60_rst0,
    input [C_INPUT_BRAM_60_WIDTH/8-1:0] ap_bram_iarg_60_we0,
    input ap_bram_iarg_60_en0,
    input [C_INPUT_BRAM_60_ADDR_WIDTH-1:0] ap_bram_iarg_60_addr1,
    input [C_INPUT_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_din1,
    output [C_INPUT_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_dout1,
    input ap_bram_iarg_60_clk1,
    input ap_bram_iarg_60_rst1,
    input [C_INPUT_BRAM_60_WIDTH/8-1:0] ap_bram_iarg_60_we1,
    input ap_bram_iarg_60_en1,
    //input AXI-Stream to BRAM interface 61
    input s_axis_bram_61_tlast,
    input s_axis_bram_61_tvalid,
    input [C_INPUT_BRAM_61_DMWIDTH/8-1:0] s_axis_bram_61_tkeep,
    input [C_INPUT_BRAM_61_DMWIDTH/8-1:0] s_axis_bram_61_tstrb,
    input [C_INPUT_BRAM_61_DMWIDTH-1:0] s_axis_bram_61_tdata,
    output s_axis_bram_61_tready,
    input [C_INPUT_BRAM_61_ADDR_WIDTH-1:0] ap_bram_iarg_61_addr0,
    input [C_INPUT_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_din0,
    output [C_INPUT_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_dout0,
    input ap_bram_iarg_61_clk0,
    input ap_bram_iarg_61_rst0,
    input [C_INPUT_BRAM_61_WIDTH/8-1:0] ap_bram_iarg_61_we0,
    input ap_bram_iarg_61_en0,
    input [C_INPUT_BRAM_61_ADDR_WIDTH-1:0] ap_bram_iarg_61_addr1,
    input [C_INPUT_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_din1,
    output [C_INPUT_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_dout1,
    input ap_bram_iarg_61_clk1,
    input ap_bram_iarg_61_rst1,
    input [C_INPUT_BRAM_61_WIDTH/8-1:0] ap_bram_iarg_61_we1,
    input ap_bram_iarg_61_en1,
    //input AXI-Stream to BRAM interface 62
    input s_axis_bram_62_tlast,
    input s_axis_bram_62_tvalid,
    input [C_INPUT_BRAM_62_DMWIDTH/8-1:0] s_axis_bram_62_tkeep,
    input [C_INPUT_BRAM_62_DMWIDTH/8-1:0] s_axis_bram_62_tstrb,
    input [C_INPUT_BRAM_62_DMWIDTH-1:0] s_axis_bram_62_tdata,
    output s_axis_bram_62_tready,
    input [C_INPUT_BRAM_62_ADDR_WIDTH-1:0] ap_bram_iarg_62_addr0,
    input [C_INPUT_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_din0,
    output [C_INPUT_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_dout0,
    input ap_bram_iarg_62_clk0,
    input ap_bram_iarg_62_rst0,
    input [C_INPUT_BRAM_62_WIDTH/8-1:0] ap_bram_iarg_62_we0,
    input ap_bram_iarg_62_en0,
    input [C_INPUT_BRAM_62_ADDR_WIDTH-1:0] ap_bram_iarg_62_addr1,
    input [C_INPUT_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_din1,
    output [C_INPUT_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_dout1,
    input ap_bram_iarg_62_clk1,
    input ap_bram_iarg_62_rst1,
    input [C_INPUT_BRAM_62_WIDTH/8-1:0] ap_bram_iarg_62_we1,
    input ap_bram_iarg_62_en1,
    //input AXI-Stream to BRAM interface 63
    input s_axis_bram_63_tlast,
    input s_axis_bram_63_tvalid,
    input [C_INPUT_BRAM_63_DMWIDTH/8-1:0] s_axis_bram_63_tkeep,
    input [C_INPUT_BRAM_63_DMWIDTH/8-1:0] s_axis_bram_63_tstrb,
    input [C_INPUT_BRAM_63_DMWIDTH-1:0] s_axis_bram_63_tdata,
    output s_axis_bram_63_tready,
    input [C_INPUT_BRAM_63_ADDR_WIDTH-1:0] ap_bram_iarg_63_addr0,
    input [C_INPUT_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_din0,
    output [C_INPUT_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_dout0,
    input ap_bram_iarg_63_clk0,
    input ap_bram_iarg_63_rst0,
    input [C_INPUT_BRAM_63_WIDTH/8-1:0] ap_bram_iarg_63_we0,
    input ap_bram_iarg_63_en0,
    input [C_INPUT_BRAM_63_ADDR_WIDTH-1:0] ap_bram_iarg_63_addr1,
    input [C_INPUT_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_din1,
    output [C_INPUT_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_dout1,
    input ap_bram_iarg_63_clk1,
    input ap_bram_iarg_63_rst1,
    input [C_INPUT_BRAM_63_WIDTH/8-1:0] ap_bram_iarg_63_we1,
    input ap_bram_iarg_63_en1,
    //input AXI-Stream to BRAM interface 64
    input s_axis_bram_64_tlast,
    input s_axis_bram_64_tvalid,
    input [C_INPUT_BRAM_64_DMWIDTH/8-1:0] s_axis_bram_64_tkeep,
    input [C_INPUT_BRAM_64_DMWIDTH/8-1:0] s_axis_bram_64_tstrb,
    input [C_INPUT_BRAM_64_DMWIDTH-1:0] s_axis_bram_64_tdata,
    output s_axis_bram_64_tready,
    input [C_INPUT_BRAM_64_ADDR_WIDTH-1:0] ap_bram_iarg_64_addr0,
    input [C_INPUT_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_din0,
    output [C_INPUT_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_dout0,
    input ap_bram_iarg_64_clk0,
    input ap_bram_iarg_64_rst0,
    input [C_INPUT_BRAM_64_WIDTH/8-1:0] ap_bram_iarg_64_we0,
    input ap_bram_iarg_64_en0,
    input [C_INPUT_BRAM_64_ADDR_WIDTH-1:0] ap_bram_iarg_64_addr1,
    input [C_INPUT_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_din1,
    output [C_INPUT_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_dout1,
    input ap_bram_iarg_64_clk1,
    input ap_bram_iarg_64_rst1,
    input [C_INPUT_BRAM_64_WIDTH/8-1:0] ap_bram_iarg_64_we1,
    input ap_bram_iarg_64_en1,
    //input AXI-Stream to BRAM interface 65
    input s_axis_bram_65_tlast,
    input s_axis_bram_65_tvalid,
    input [C_INPUT_BRAM_65_DMWIDTH/8-1:0] s_axis_bram_65_tkeep,
    input [C_INPUT_BRAM_65_DMWIDTH/8-1:0] s_axis_bram_65_tstrb,
    input [C_INPUT_BRAM_65_DMWIDTH-1:0] s_axis_bram_65_tdata,
    output s_axis_bram_65_tready,
    input [C_INPUT_BRAM_65_ADDR_WIDTH-1:0] ap_bram_iarg_65_addr0,
    input [C_INPUT_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_din0,
    output [C_INPUT_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_dout0,
    input ap_bram_iarg_65_clk0,
    input ap_bram_iarg_65_rst0,
    input [C_INPUT_BRAM_65_WIDTH/8-1:0] ap_bram_iarg_65_we0,
    input ap_bram_iarg_65_en0,
    input [C_INPUT_BRAM_65_ADDR_WIDTH-1:0] ap_bram_iarg_65_addr1,
    input [C_INPUT_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_din1,
    output [C_INPUT_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_dout1,
    input ap_bram_iarg_65_clk1,
    input ap_bram_iarg_65_rst1,
    input [C_INPUT_BRAM_65_WIDTH/8-1:0] ap_bram_iarg_65_we1,
    input ap_bram_iarg_65_en1,
    //input AXI-Stream to BRAM interface 66
    input s_axis_bram_66_tlast,
    input s_axis_bram_66_tvalid,
    input [C_INPUT_BRAM_66_DMWIDTH/8-1:0] s_axis_bram_66_tkeep,
    input [C_INPUT_BRAM_66_DMWIDTH/8-1:0] s_axis_bram_66_tstrb,
    input [C_INPUT_BRAM_66_DMWIDTH-1:0] s_axis_bram_66_tdata,
    output s_axis_bram_66_tready,
    input [C_INPUT_BRAM_66_ADDR_WIDTH-1:0] ap_bram_iarg_66_addr0,
    input [C_INPUT_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_din0,
    output [C_INPUT_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_dout0,
    input ap_bram_iarg_66_clk0,
    input ap_bram_iarg_66_rst0,
    input [C_INPUT_BRAM_66_WIDTH/8-1:0] ap_bram_iarg_66_we0,
    input ap_bram_iarg_66_en0,
    input [C_INPUT_BRAM_66_ADDR_WIDTH-1:0] ap_bram_iarg_66_addr1,
    input [C_INPUT_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_din1,
    output [C_INPUT_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_dout1,
    input ap_bram_iarg_66_clk1,
    input ap_bram_iarg_66_rst1,
    input [C_INPUT_BRAM_66_WIDTH/8-1:0] ap_bram_iarg_66_we1,
    input ap_bram_iarg_66_en1,
    //input AXI-Stream to BRAM interface 67
    input s_axis_bram_67_tlast,
    input s_axis_bram_67_tvalid,
    input [C_INPUT_BRAM_67_DMWIDTH/8-1:0] s_axis_bram_67_tkeep,
    input [C_INPUT_BRAM_67_DMWIDTH/8-1:0] s_axis_bram_67_tstrb,
    input [C_INPUT_BRAM_67_DMWIDTH-1:0] s_axis_bram_67_tdata,
    output s_axis_bram_67_tready,
    input [C_INPUT_BRAM_67_ADDR_WIDTH-1:0] ap_bram_iarg_67_addr0,
    input [C_INPUT_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_din0,
    output [C_INPUT_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_dout0,
    input ap_bram_iarg_67_clk0,
    input ap_bram_iarg_67_rst0,
    input [C_INPUT_BRAM_67_WIDTH/8-1:0] ap_bram_iarg_67_we0,
    input ap_bram_iarg_67_en0,
    input [C_INPUT_BRAM_67_ADDR_WIDTH-1:0] ap_bram_iarg_67_addr1,
    input [C_INPUT_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_din1,
    output [C_INPUT_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_dout1,
    input ap_bram_iarg_67_clk1,
    input ap_bram_iarg_67_rst1,
    input [C_INPUT_BRAM_67_WIDTH/8-1:0] ap_bram_iarg_67_we1,
    input ap_bram_iarg_67_en1,
    //input AXI-Stream to BRAM interface 68
    input s_axis_bram_68_tlast,
    input s_axis_bram_68_tvalid,
    input [C_INPUT_BRAM_68_DMWIDTH/8-1:0] s_axis_bram_68_tkeep,
    input [C_INPUT_BRAM_68_DMWIDTH/8-1:0] s_axis_bram_68_tstrb,
    input [C_INPUT_BRAM_68_DMWIDTH-1:0] s_axis_bram_68_tdata,
    output s_axis_bram_68_tready,
    input [C_INPUT_BRAM_68_ADDR_WIDTH-1:0] ap_bram_iarg_68_addr0,
    input [C_INPUT_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_din0,
    output [C_INPUT_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_dout0,
    input ap_bram_iarg_68_clk0,
    input ap_bram_iarg_68_rst0,
    input [C_INPUT_BRAM_68_WIDTH/8-1:0] ap_bram_iarg_68_we0,
    input ap_bram_iarg_68_en0,
    input [C_INPUT_BRAM_68_ADDR_WIDTH-1:0] ap_bram_iarg_68_addr1,
    input [C_INPUT_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_din1,
    output [C_INPUT_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_dout1,
    input ap_bram_iarg_68_clk1,
    input ap_bram_iarg_68_rst1,
    input [C_INPUT_BRAM_68_WIDTH/8-1:0] ap_bram_iarg_68_we1,
    input ap_bram_iarg_68_en1,
    //input AXI-Stream to BRAM interface 69
    input s_axis_bram_69_tlast,
    input s_axis_bram_69_tvalid,
    input [C_INPUT_BRAM_69_DMWIDTH/8-1:0] s_axis_bram_69_tkeep,
    input [C_INPUT_BRAM_69_DMWIDTH/8-1:0] s_axis_bram_69_tstrb,
    input [C_INPUT_BRAM_69_DMWIDTH-1:0] s_axis_bram_69_tdata,
    output s_axis_bram_69_tready,
    input [C_INPUT_BRAM_69_ADDR_WIDTH-1:0] ap_bram_iarg_69_addr0,
    input [C_INPUT_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_din0,
    output [C_INPUT_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_dout0,
    input ap_bram_iarg_69_clk0,
    input ap_bram_iarg_69_rst0,
    input [C_INPUT_BRAM_69_WIDTH/8-1:0] ap_bram_iarg_69_we0,
    input ap_bram_iarg_69_en0,
    input [C_INPUT_BRAM_69_ADDR_WIDTH-1:0] ap_bram_iarg_69_addr1,
    input [C_INPUT_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_din1,
    output [C_INPUT_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_dout1,
    input ap_bram_iarg_69_clk1,
    input ap_bram_iarg_69_rst1,
    input [C_INPUT_BRAM_69_WIDTH/8-1:0] ap_bram_iarg_69_we1,
    input ap_bram_iarg_69_en1,
    //input AXI-Stream to BRAM interface 70
    input s_axis_bram_70_tlast,
    input s_axis_bram_70_tvalid,
    input [C_INPUT_BRAM_70_DMWIDTH/8-1:0] s_axis_bram_70_tkeep,
    input [C_INPUT_BRAM_70_DMWIDTH/8-1:0] s_axis_bram_70_tstrb,
    input [C_INPUT_BRAM_70_DMWIDTH-1:0] s_axis_bram_70_tdata,
    output s_axis_bram_70_tready,
    input [C_INPUT_BRAM_70_ADDR_WIDTH-1:0] ap_bram_iarg_70_addr0,
    input [C_INPUT_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_din0,
    output [C_INPUT_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_dout0,
    input ap_bram_iarg_70_clk0,
    input ap_bram_iarg_70_rst0,
    input [C_INPUT_BRAM_70_WIDTH/8-1:0] ap_bram_iarg_70_we0,
    input ap_bram_iarg_70_en0,
    input [C_INPUT_BRAM_70_ADDR_WIDTH-1:0] ap_bram_iarg_70_addr1,
    input [C_INPUT_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_din1,
    output [C_INPUT_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_dout1,
    input ap_bram_iarg_70_clk1,
    input ap_bram_iarg_70_rst1,
    input [C_INPUT_BRAM_70_WIDTH/8-1:0] ap_bram_iarg_70_we1,
    input ap_bram_iarg_70_en1,
    //input AXI-Stream to BRAM interface 71
    input s_axis_bram_71_tlast,
    input s_axis_bram_71_tvalid,
    input [C_INPUT_BRAM_71_DMWIDTH/8-1:0] s_axis_bram_71_tkeep,
    input [C_INPUT_BRAM_71_DMWIDTH/8-1:0] s_axis_bram_71_tstrb,
    input [C_INPUT_BRAM_71_DMWIDTH-1:0] s_axis_bram_71_tdata,
    output s_axis_bram_71_tready,
    input [C_INPUT_BRAM_71_ADDR_WIDTH-1:0] ap_bram_iarg_71_addr0,
    input [C_INPUT_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_din0,
    output [C_INPUT_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_dout0,
    input ap_bram_iarg_71_clk0,
    input ap_bram_iarg_71_rst0,
    input [C_INPUT_BRAM_71_WIDTH/8-1:0] ap_bram_iarg_71_we0,
    input ap_bram_iarg_71_en0,
    input [C_INPUT_BRAM_71_ADDR_WIDTH-1:0] ap_bram_iarg_71_addr1,
    input [C_INPUT_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_din1,
    output [C_INPUT_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_dout1,
    input ap_bram_iarg_71_clk1,
    input ap_bram_iarg_71_rst1,
    input [C_INPUT_BRAM_71_WIDTH/8-1:0] ap_bram_iarg_71_we1,
    input ap_bram_iarg_71_en1,
    //input AXI-Stream to BRAM interface 72
    input s_axis_bram_72_tlast,
    input s_axis_bram_72_tvalid,
    input [C_INPUT_BRAM_72_DMWIDTH/8-1:0] s_axis_bram_72_tkeep,
    input [C_INPUT_BRAM_72_DMWIDTH/8-1:0] s_axis_bram_72_tstrb,
    input [C_INPUT_BRAM_72_DMWIDTH-1:0] s_axis_bram_72_tdata,
    output s_axis_bram_72_tready,
    input [C_INPUT_BRAM_72_ADDR_WIDTH-1:0] ap_bram_iarg_72_addr0,
    input [C_INPUT_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_din0,
    output [C_INPUT_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_dout0,
    input ap_bram_iarg_72_clk0,
    input ap_bram_iarg_72_rst0,
    input [C_INPUT_BRAM_72_WIDTH/8-1:0] ap_bram_iarg_72_we0,
    input ap_bram_iarg_72_en0,
    input [C_INPUT_BRAM_72_ADDR_WIDTH-1:0] ap_bram_iarg_72_addr1,
    input [C_INPUT_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_din1,
    output [C_INPUT_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_dout1,
    input ap_bram_iarg_72_clk1,
    input ap_bram_iarg_72_rst1,
    input [C_INPUT_BRAM_72_WIDTH/8-1:0] ap_bram_iarg_72_we1,
    input ap_bram_iarg_72_en1,
    //input AXI-Stream to BRAM interface 73
    input s_axis_bram_73_tlast,
    input s_axis_bram_73_tvalid,
    input [C_INPUT_BRAM_73_DMWIDTH/8-1:0] s_axis_bram_73_tkeep,
    input [C_INPUT_BRAM_73_DMWIDTH/8-1:0] s_axis_bram_73_tstrb,
    input [C_INPUT_BRAM_73_DMWIDTH-1:0] s_axis_bram_73_tdata,
    output s_axis_bram_73_tready,
    input [C_INPUT_BRAM_73_ADDR_WIDTH-1:0] ap_bram_iarg_73_addr0,
    input [C_INPUT_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_din0,
    output [C_INPUT_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_dout0,
    input ap_bram_iarg_73_clk0,
    input ap_bram_iarg_73_rst0,
    input [C_INPUT_BRAM_73_WIDTH/8-1:0] ap_bram_iarg_73_we0,
    input ap_bram_iarg_73_en0,
    input [C_INPUT_BRAM_73_ADDR_WIDTH-1:0] ap_bram_iarg_73_addr1,
    input [C_INPUT_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_din1,
    output [C_INPUT_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_dout1,
    input ap_bram_iarg_73_clk1,
    input ap_bram_iarg_73_rst1,
    input [C_INPUT_BRAM_73_WIDTH/8-1:0] ap_bram_iarg_73_we1,
    input ap_bram_iarg_73_en1,
    //input AXI-Stream to BRAM interface 74
    input s_axis_bram_74_tlast,
    input s_axis_bram_74_tvalid,
    input [C_INPUT_BRAM_74_DMWIDTH/8-1:0] s_axis_bram_74_tkeep,
    input [C_INPUT_BRAM_74_DMWIDTH/8-1:0] s_axis_bram_74_tstrb,
    input [C_INPUT_BRAM_74_DMWIDTH-1:0] s_axis_bram_74_tdata,
    output s_axis_bram_74_tready,
    input [C_INPUT_BRAM_74_ADDR_WIDTH-1:0] ap_bram_iarg_74_addr0,
    input [C_INPUT_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_din0,
    output [C_INPUT_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_dout0,
    input ap_bram_iarg_74_clk0,
    input ap_bram_iarg_74_rst0,
    input [C_INPUT_BRAM_74_WIDTH/8-1:0] ap_bram_iarg_74_we0,
    input ap_bram_iarg_74_en0,
    input [C_INPUT_BRAM_74_ADDR_WIDTH-1:0] ap_bram_iarg_74_addr1,
    input [C_INPUT_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_din1,
    output [C_INPUT_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_dout1,
    input ap_bram_iarg_74_clk1,
    input ap_bram_iarg_74_rst1,
    input [C_INPUT_BRAM_74_WIDTH/8-1:0] ap_bram_iarg_74_we1,
    input ap_bram_iarg_74_en1,
    //input AXI-Stream to BRAM interface 75
    input s_axis_bram_75_tlast,
    input s_axis_bram_75_tvalid,
    input [C_INPUT_BRAM_75_DMWIDTH/8-1:0] s_axis_bram_75_tkeep,
    input [C_INPUT_BRAM_75_DMWIDTH/8-1:0] s_axis_bram_75_tstrb,
    input [C_INPUT_BRAM_75_DMWIDTH-1:0] s_axis_bram_75_tdata,
    output s_axis_bram_75_tready,
    input [C_INPUT_BRAM_75_ADDR_WIDTH-1:0] ap_bram_iarg_75_addr0,
    input [C_INPUT_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_din0,
    output [C_INPUT_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_dout0,
    input ap_bram_iarg_75_clk0,
    input ap_bram_iarg_75_rst0,
    input [C_INPUT_BRAM_75_WIDTH/8-1:0] ap_bram_iarg_75_we0,
    input ap_bram_iarg_75_en0,
    input [C_INPUT_BRAM_75_ADDR_WIDTH-1:0] ap_bram_iarg_75_addr1,
    input [C_INPUT_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_din1,
    output [C_INPUT_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_dout1,
    input ap_bram_iarg_75_clk1,
    input ap_bram_iarg_75_rst1,
    input [C_INPUT_BRAM_75_WIDTH/8-1:0] ap_bram_iarg_75_we1,
    input ap_bram_iarg_75_en1,
    //input AXI-Stream to BRAM interface 76
    input s_axis_bram_76_tlast,
    input s_axis_bram_76_tvalid,
    input [C_INPUT_BRAM_76_DMWIDTH/8-1:0] s_axis_bram_76_tkeep,
    input [C_INPUT_BRAM_76_DMWIDTH/8-1:0] s_axis_bram_76_tstrb,
    input [C_INPUT_BRAM_76_DMWIDTH-1:0] s_axis_bram_76_tdata,
    output s_axis_bram_76_tready,
    input [C_INPUT_BRAM_76_ADDR_WIDTH-1:0] ap_bram_iarg_76_addr0,
    input [C_INPUT_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_din0,
    output [C_INPUT_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_dout0,
    input ap_bram_iarg_76_clk0,
    input ap_bram_iarg_76_rst0,
    input [C_INPUT_BRAM_76_WIDTH/8-1:0] ap_bram_iarg_76_we0,
    input ap_bram_iarg_76_en0,
    input [C_INPUT_BRAM_76_ADDR_WIDTH-1:0] ap_bram_iarg_76_addr1,
    input [C_INPUT_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_din1,
    output [C_INPUT_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_dout1,
    input ap_bram_iarg_76_clk1,
    input ap_bram_iarg_76_rst1,
    input [C_INPUT_BRAM_76_WIDTH/8-1:0] ap_bram_iarg_76_we1,
    input ap_bram_iarg_76_en1,
    //input AXI-Stream to BRAM interface 77
    input s_axis_bram_77_tlast,
    input s_axis_bram_77_tvalid,
    input [C_INPUT_BRAM_77_DMWIDTH/8-1:0] s_axis_bram_77_tkeep,
    input [C_INPUT_BRAM_77_DMWIDTH/8-1:0] s_axis_bram_77_tstrb,
    input [C_INPUT_BRAM_77_DMWIDTH-1:0] s_axis_bram_77_tdata,
    output s_axis_bram_77_tready,
    input [C_INPUT_BRAM_77_ADDR_WIDTH-1:0] ap_bram_iarg_77_addr0,
    input [C_INPUT_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_din0,
    output [C_INPUT_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_dout0,
    input ap_bram_iarg_77_clk0,
    input ap_bram_iarg_77_rst0,
    input [C_INPUT_BRAM_77_WIDTH/8-1:0] ap_bram_iarg_77_we0,
    input ap_bram_iarg_77_en0,
    input [C_INPUT_BRAM_77_ADDR_WIDTH-1:0] ap_bram_iarg_77_addr1,
    input [C_INPUT_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_din1,
    output [C_INPUT_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_dout1,
    input ap_bram_iarg_77_clk1,
    input ap_bram_iarg_77_rst1,
    input [C_INPUT_BRAM_77_WIDTH/8-1:0] ap_bram_iarg_77_we1,
    input ap_bram_iarg_77_en1,
    //input AXI-Stream to BRAM interface 78
    input s_axis_bram_78_tlast,
    input s_axis_bram_78_tvalid,
    input [C_INPUT_BRAM_78_DMWIDTH/8-1:0] s_axis_bram_78_tkeep,
    input [C_INPUT_BRAM_78_DMWIDTH/8-1:0] s_axis_bram_78_tstrb,
    input [C_INPUT_BRAM_78_DMWIDTH-1:0] s_axis_bram_78_tdata,
    output s_axis_bram_78_tready,
    input [C_INPUT_BRAM_78_ADDR_WIDTH-1:0] ap_bram_iarg_78_addr0,
    input [C_INPUT_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_din0,
    output [C_INPUT_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_dout0,
    input ap_bram_iarg_78_clk0,
    input ap_bram_iarg_78_rst0,
    input [C_INPUT_BRAM_78_WIDTH/8-1:0] ap_bram_iarg_78_we0,
    input ap_bram_iarg_78_en0,
    input [C_INPUT_BRAM_78_ADDR_WIDTH-1:0] ap_bram_iarg_78_addr1,
    input [C_INPUT_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_din1,
    output [C_INPUT_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_dout1,
    input ap_bram_iarg_78_clk1,
    input ap_bram_iarg_78_rst1,
    input [C_INPUT_BRAM_78_WIDTH/8-1:0] ap_bram_iarg_78_we1,
    input ap_bram_iarg_78_en1,
    //input AXI-Stream to BRAM interface 79
    input s_axis_bram_79_tlast,
    input s_axis_bram_79_tvalid,
    input [C_INPUT_BRAM_79_DMWIDTH/8-1:0] s_axis_bram_79_tkeep,
    input [C_INPUT_BRAM_79_DMWIDTH/8-1:0] s_axis_bram_79_tstrb,
    input [C_INPUT_BRAM_79_DMWIDTH-1:0] s_axis_bram_79_tdata,
    output s_axis_bram_79_tready,
    input [C_INPUT_BRAM_79_ADDR_WIDTH-1:0] ap_bram_iarg_79_addr0,
    input [C_INPUT_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_din0,
    output [C_INPUT_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_dout0,
    input ap_bram_iarg_79_clk0,
    input ap_bram_iarg_79_rst0,
    input [C_INPUT_BRAM_79_WIDTH/8-1:0] ap_bram_iarg_79_we0,
    input ap_bram_iarg_79_en0,
    input [C_INPUT_BRAM_79_ADDR_WIDTH-1:0] ap_bram_iarg_79_addr1,
    input [C_INPUT_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_din1,
    output [C_INPUT_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_dout1,
    input ap_bram_iarg_79_clk1,
    input ap_bram_iarg_79_rst1,
    input [C_INPUT_BRAM_79_WIDTH/8-1:0] ap_bram_iarg_79_we1,
    input ap_bram_iarg_79_en1,
    //input AXI-Stream to BRAM interface 80
    input s_axis_bram_80_tlast,
    input s_axis_bram_80_tvalid,
    input [C_INPUT_BRAM_80_DMWIDTH/8-1:0] s_axis_bram_80_tkeep,
    input [C_INPUT_BRAM_80_DMWIDTH/8-1:0] s_axis_bram_80_tstrb,
    input [C_INPUT_BRAM_80_DMWIDTH-1:0] s_axis_bram_80_tdata,
    output s_axis_bram_80_tready,
    input [C_INPUT_BRAM_80_ADDR_WIDTH-1:0] ap_bram_iarg_80_addr0,
    input [C_INPUT_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_din0,
    output [C_INPUT_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_dout0,
    input ap_bram_iarg_80_clk0,
    input ap_bram_iarg_80_rst0,
    input [C_INPUT_BRAM_80_WIDTH/8-1:0] ap_bram_iarg_80_we0,
    input ap_bram_iarg_80_en0,
    input [C_INPUT_BRAM_80_ADDR_WIDTH-1:0] ap_bram_iarg_80_addr1,
    input [C_INPUT_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_din1,
    output [C_INPUT_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_dout1,
    input ap_bram_iarg_80_clk1,
    input ap_bram_iarg_80_rst1,
    input [C_INPUT_BRAM_80_WIDTH/8-1:0] ap_bram_iarg_80_we1,
    input ap_bram_iarg_80_en1,
    //input AXI-Stream to BRAM interface 81
    input s_axis_bram_81_tlast,
    input s_axis_bram_81_tvalid,
    input [C_INPUT_BRAM_81_DMWIDTH/8-1:0] s_axis_bram_81_tkeep,
    input [C_INPUT_BRAM_81_DMWIDTH/8-1:0] s_axis_bram_81_tstrb,
    input [C_INPUT_BRAM_81_DMWIDTH-1:0] s_axis_bram_81_tdata,
    output s_axis_bram_81_tready,
    input [C_INPUT_BRAM_81_ADDR_WIDTH-1:0] ap_bram_iarg_81_addr0,
    input [C_INPUT_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_din0,
    output [C_INPUT_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_dout0,
    input ap_bram_iarg_81_clk0,
    input ap_bram_iarg_81_rst0,
    input [C_INPUT_BRAM_81_WIDTH/8-1:0] ap_bram_iarg_81_we0,
    input ap_bram_iarg_81_en0,
    input [C_INPUT_BRAM_81_ADDR_WIDTH-1:0] ap_bram_iarg_81_addr1,
    input [C_INPUT_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_din1,
    output [C_INPUT_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_dout1,
    input ap_bram_iarg_81_clk1,
    input ap_bram_iarg_81_rst1,
    input [C_INPUT_BRAM_81_WIDTH/8-1:0] ap_bram_iarg_81_we1,
    input ap_bram_iarg_81_en1,
    //input AXI-Stream to BRAM interface 82
    input s_axis_bram_82_tlast,
    input s_axis_bram_82_tvalid,
    input [C_INPUT_BRAM_82_DMWIDTH/8-1:0] s_axis_bram_82_tkeep,
    input [C_INPUT_BRAM_82_DMWIDTH/8-1:0] s_axis_bram_82_tstrb,
    input [C_INPUT_BRAM_82_DMWIDTH-1:0] s_axis_bram_82_tdata,
    output s_axis_bram_82_tready,
    input [C_INPUT_BRAM_82_ADDR_WIDTH-1:0] ap_bram_iarg_82_addr0,
    input [C_INPUT_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_din0,
    output [C_INPUT_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_dout0,
    input ap_bram_iarg_82_clk0,
    input ap_bram_iarg_82_rst0,
    input [C_INPUT_BRAM_82_WIDTH/8-1:0] ap_bram_iarg_82_we0,
    input ap_bram_iarg_82_en0,
    input [C_INPUT_BRAM_82_ADDR_WIDTH-1:0] ap_bram_iarg_82_addr1,
    input [C_INPUT_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_din1,
    output [C_INPUT_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_dout1,
    input ap_bram_iarg_82_clk1,
    input ap_bram_iarg_82_rst1,
    input [C_INPUT_BRAM_82_WIDTH/8-1:0] ap_bram_iarg_82_we1,
    input ap_bram_iarg_82_en1,
    //input AXI-Stream to BRAM interface 83
    input s_axis_bram_83_tlast,
    input s_axis_bram_83_tvalid,
    input [C_INPUT_BRAM_83_DMWIDTH/8-1:0] s_axis_bram_83_tkeep,
    input [C_INPUT_BRAM_83_DMWIDTH/8-1:0] s_axis_bram_83_tstrb,
    input [C_INPUT_BRAM_83_DMWIDTH-1:0] s_axis_bram_83_tdata,
    output s_axis_bram_83_tready,
    input [C_INPUT_BRAM_83_ADDR_WIDTH-1:0] ap_bram_iarg_83_addr0,
    input [C_INPUT_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_din0,
    output [C_INPUT_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_dout0,
    input ap_bram_iarg_83_clk0,
    input ap_bram_iarg_83_rst0,
    input [C_INPUT_BRAM_83_WIDTH/8-1:0] ap_bram_iarg_83_we0,
    input ap_bram_iarg_83_en0,
    input [C_INPUT_BRAM_83_ADDR_WIDTH-1:0] ap_bram_iarg_83_addr1,
    input [C_INPUT_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_din1,
    output [C_INPUT_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_dout1,
    input ap_bram_iarg_83_clk1,
    input ap_bram_iarg_83_rst1,
    input [C_INPUT_BRAM_83_WIDTH/8-1:0] ap_bram_iarg_83_we1,
    input ap_bram_iarg_83_en1,
    //input AXI-Stream to BRAM interface 84
    input s_axis_bram_84_tlast,
    input s_axis_bram_84_tvalid,
    input [C_INPUT_BRAM_84_DMWIDTH/8-1:0] s_axis_bram_84_tkeep,
    input [C_INPUT_BRAM_84_DMWIDTH/8-1:0] s_axis_bram_84_tstrb,
    input [C_INPUT_BRAM_84_DMWIDTH-1:0] s_axis_bram_84_tdata,
    output s_axis_bram_84_tready,
    input [C_INPUT_BRAM_84_ADDR_WIDTH-1:0] ap_bram_iarg_84_addr0,
    input [C_INPUT_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_din0,
    output [C_INPUT_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_dout0,
    input ap_bram_iarg_84_clk0,
    input ap_bram_iarg_84_rst0,
    input [C_INPUT_BRAM_84_WIDTH/8-1:0] ap_bram_iarg_84_we0,
    input ap_bram_iarg_84_en0,
    input [C_INPUT_BRAM_84_ADDR_WIDTH-1:0] ap_bram_iarg_84_addr1,
    input [C_INPUT_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_din1,
    output [C_INPUT_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_dout1,
    input ap_bram_iarg_84_clk1,
    input ap_bram_iarg_84_rst1,
    input [C_INPUT_BRAM_84_WIDTH/8-1:0] ap_bram_iarg_84_we1,
    input ap_bram_iarg_84_en1,
    //input AXI-Stream to BRAM interface 85
    input s_axis_bram_85_tlast,
    input s_axis_bram_85_tvalid,
    input [C_INPUT_BRAM_85_DMWIDTH/8-1:0] s_axis_bram_85_tkeep,
    input [C_INPUT_BRAM_85_DMWIDTH/8-1:0] s_axis_bram_85_tstrb,
    input [C_INPUT_BRAM_85_DMWIDTH-1:0] s_axis_bram_85_tdata,
    output s_axis_bram_85_tready,
    input [C_INPUT_BRAM_85_ADDR_WIDTH-1:0] ap_bram_iarg_85_addr0,
    input [C_INPUT_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_din0,
    output [C_INPUT_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_dout0,
    input ap_bram_iarg_85_clk0,
    input ap_bram_iarg_85_rst0,
    input [C_INPUT_BRAM_85_WIDTH/8-1:0] ap_bram_iarg_85_we0,
    input ap_bram_iarg_85_en0,
    input [C_INPUT_BRAM_85_ADDR_WIDTH-1:0] ap_bram_iarg_85_addr1,
    input [C_INPUT_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_din1,
    output [C_INPUT_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_dout1,
    input ap_bram_iarg_85_clk1,
    input ap_bram_iarg_85_rst1,
    input [C_INPUT_BRAM_85_WIDTH/8-1:0] ap_bram_iarg_85_we1,
    input ap_bram_iarg_85_en1,
    //input AXI-Stream to BRAM interface 86
    input s_axis_bram_86_tlast,
    input s_axis_bram_86_tvalid,
    input [C_INPUT_BRAM_86_DMWIDTH/8-1:0] s_axis_bram_86_tkeep,
    input [C_INPUT_BRAM_86_DMWIDTH/8-1:0] s_axis_bram_86_tstrb,
    input [C_INPUT_BRAM_86_DMWIDTH-1:0] s_axis_bram_86_tdata,
    output s_axis_bram_86_tready,
    input [C_INPUT_BRAM_86_ADDR_WIDTH-1:0] ap_bram_iarg_86_addr0,
    input [C_INPUT_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_din0,
    output [C_INPUT_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_dout0,
    input ap_bram_iarg_86_clk0,
    input ap_bram_iarg_86_rst0,
    input [C_INPUT_BRAM_86_WIDTH/8-1:0] ap_bram_iarg_86_we0,
    input ap_bram_iarg_86_en0,
    input [C_INPUT_BRAM_86_ADDR_WIDTH-1:0] ap_bram_iarg_86_addr1,
    input [C_INPUT_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_din1,
    output [C_INPUT_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_dout1,
    input ap_bram_iarg_86_clk1,
    input ap_bram_iarg_86_rst1,
    input [C_INPUT_BRAM_86_WIDTH/8-1:0] ap_bram_iarg_86_we1,
    input ap_bram_iarg_86_en1,
    //input AXI-Stream to BRAM interface 87
    input s_axis_bram_87_tlast,
    input s_axis_bram_87_tvalid,
    input [C_INPUT_BRAM_87_DMWIDTH/8-1:0] s_axis_bram_87_tkeep,
    input [C_INPUT_BRAM_87_DMWIDTH/8-1:0] s_axis_bram_87_tstrb,
    input [C_INPUT_BRAM_87_DMWIDTH-1:0] s_axis_bram_87_tdata,
    output s_axis_bram_87_tready,
    input [C_INPUT_BRAM_87_ADDR_WIDTH-1:0] ap_bram_iarg_87_addr0,
    input [C_INPUT_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_din0,
    output [C_INPUT_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_dout0,
    input ap_bram_iarg_87_clk0,
    input ap_bram_iarg_87_rst0,
    input [C_INPUT_BRAM_87_WIDTH/8-1:0] ap_bram_iarg_87_we0,
    input ap_bram_iarg_87_en0,
    input [C_INPUT_BRAM_87_ADDR_WIDTH-1:0] ap_bram_iarg_87_addr1,
    input [C_INPUT_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_din1,
    output [C_INPUT_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_dout1,
    input ap_bram_iarg_87_clk1,
    input ap_bram_iarg_87_rst1,
    input [C_INPUT_BRAM_87_WIDTH/8-1:0] ap_bram_iarg_87_we1,
    input ap_bram_iarg_87_en1,
    //input AXI-Stream to BRAM interface 88
    input s_axis_bram_88_tlast,
    input s_axis_bram_88_tvalid,
    input [C_INPUT_BRAM_88_DMWIDTH/8-1:0] s_axis_bram_88_tkeep,
    input [C_INPUT_BRAM_88_DMWIDTH/8-1:0] s_axis_bram_88_tstrb,
    input [C_INPUT_BRAM_88_DMWIDTH-1:0] s_axis_bram_88_tdata,
    output s_axis_bram_88_tready,
    input [C_INPUT_BRAM_88_ADDR_WIDTH-1:0] ap_bram_iarg_88_addr0,
    input [C_INPUT_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_din0,
    output [C_INPUT_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_dout0,
    input ap_bram_iarg_88_clk0,
    input ap_bram_iarg_88_rst0,
    input [C_INPUT_BRAM_88_WIDTH/8-1:0] ap_bram_iarg_88_we0,
    input ap_bram_iarg_88_en0,
    input [C_INPUT_BRAM_88_ADDR_WIDTH-1:0] ap_bram_iarg_88_addr1,
    input [C_INPUT_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_din1,
    output [C_INPUT_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_dout1,
    input ap_bram_iarg_88_clk1,
    input ap_bram_iarg_88_rst1,
    input [C_INPUT_BRAM_88_WIDTH/8-1:0] ap_bram_iarg_88_we1,
    input ap_bram_iarg_88_en1,
    //input AXI-Stream to BRAM interface 89
    input s_axis_bram_89_tlast,
    input s_axis_bram_89_tvalid,
    input [C_INPUT_BRAM_89_DMWIDTH/8-1:0] s_axis_bram_89_tkeep,
    input [C_INPUT_BRAM_89_DMWIDTH/8-1:0] s_axis_bram_89_tstrb,
    input [C_INPUT_BRAM_89_DMWIDTH-1:0] s_axis_bram_89_tdata,
    output s_axis_bram_89_tready,
    input [C_INPUT_BRAM_89_ADDR_WIDTH-1:0] ap_bram_iarg_89_addr0,
    input [C_INPUT_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_din0,
    output [C_INPUT_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_dout0,
    input ap_bram_iarg_89_clk0,
    input ap_bram_iarg_89_rst0,
    input [C_INPUT_BRAM_89_WIDTH/8-1:0] ap_bram_iarg_89_we0,
    input ap_bram_iarg_89_en0,
    input [C_INPUT_BRAM_89_ADDR_WIDTH-1:0] ap_bram_iarg_89_addr1,
    input [C_INPUT_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_din1,
    output [C_INPUT_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_dout1,
    input ap_bram_iarg_89_clk1,
    input ap_bram_iarg_89_rst1,
    input [C_INPUT_BRAM_89_WIDTH/8-1:0] ap_bram_iarg_89_we1,
    input ap_bram_iarg_89_en1,
    //input AXI-Stream to BRAM interface 90
    input s_axis_bram_90_tlast,
    input s_axis_bram_90_tvalid,
    input [C_INPUT_BRAM_90_DMWIDTH/8-1:0] s_axis_bram_90_tkeep,
    input [C_INPUT_BRAM_90_DMWIDTH/8-1:0] s_axis_bram_90_tstrb,
    input [C_INPUT_BRAM_90_DMWIDTH-1:0] s_axis_bram_90_tdata,
    output s_axis_bram_90_tready,
    input [C_INPUT_BRAM_90_ADDR_WIDTH-1:0] ap_bram_iarg_90_addr0,
    input [C_INPUT_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_din0,
    output [C_INPUT_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_dout0,
    input ap_bram_iarg_90_clk0,
    input ap_bram_iarg_90_rst0,
    input [C_INPUT_BRAM_90_WIDTH/8-1:0] ap_bram_iarg_90_we0,
    input ap_bram_iarg_90_en0,
    input [C_INPUT_BRAM_90_ADDR_WIDTH-1:0] ap_bram_iarg_90_addr1,
    input [C_INPUT_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_din1,
    output [C_INPUT_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_dout1,
    input ap_bram_iarg_90_clk1,
    input ap_bram_iarg_90_rst1,
    input [C_INPUT_BRAM_90_WIDTH/8-1:0] ap_bram_iarg_90_we1,
    input ap_bram_iarg_90_en1,
    //input AXI-Stream to BRAM interface 91
    input s_axis_bram_91_tlast,
    input s_axis_bram_91_tvalid,
    input [C_INPUT_BRAM_91_DMWIDTH/8-1:0] s_axis_bram_91_tkeep,
    input [C_INPUT_BRAM_91_DMWIDTH/8-1:0] s_axis_bram_91_tstrb,
    input [C_INPUT_BRAM_91_DMWIDTH-1:0] s_axis_bram_91_tdata,
    output s_axis_bram_91_tready,
    input [C_INPUT_BRAM_91_ADDR_WIDTH-1:0] ap_bram_iarg_91_addr0,
    input [C_INPUT_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_din0,
    output [C_INPUT_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_dout0,
    input ap_bram_iarg_91_clk0,
    input ap_bram_iarg_91_rst0,
    input [C_INPUT_BRAM_91_WIDTH/8-1:0] ap_bram_iarg_91_we0,
    input ap_bram_iarg_91_en0,
    input [C_INPUT_BRAM_91_ADDR_WIDTH-1:0] ap_bram_iarg_91_addr1,
    input [C_INPUT_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_din1,
    output [C_INPUT_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_dout1,
    input ap_bram_iarg_91_clk1,
    input ap_bram_iarg_91_rst1,
    input [C_INPUT_BRAM_91_WIDTH/8-1:0] ap_bram_iarg_91_we1,
    input ap_bram_iarg_91_en1,
    //input AXI-Stream to BRAM interface 92
    input s_axis_bram_92_tlast,
    input s_axis_bram_92_tvalid,
    input [C_INPUT_BRAM_92_DMWIDTH/8-1:0] s_axis_bram_92_tkeep,
    input [C_INPUT_BRAM_92_DMWIDTH/8-1:0] s_axis_bram_92_tstrb,
    input [C_INPUT_BRAM_92_DMWIDTH-1:0] s_axis_bram_92_tdata,
    output s_axis_bram_92_tready,
    input [C_INPUT_BRAM_92_ADDR_WIDTH-1:0] ap_bram_iarg_92_addr0,
    input [C_INPUT_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_din0,
    output [C_INPUT_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_dout0,
    input ap_bram_iarg_92_clk0,
    input ap_bram_iarg_92_rst0,
    input [C_INPUT_BRAM_92_WIDTH/8-1:0] ap_bram_iarg_92_we0,
    input ap_bram_iarg_92_en0,
    input [C_INPUT_BRAM_92_ADDR_WIDTH-1:0] ap_bram_iarg_92_addr1,
    input [C_INPUT_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_din1,
    output [C_INPUT_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_dout1,
    input ap_bram_iarg_92_clk1,
    input ap_bram_iarg_92_rst1,
    input [C_INPUT_BRAM_92_WIDTH/8-1:0] ap_bram_iarg_92_we1,
    input ap_bram_iarg_92_en1,
    //input AXI-Stream to BRAM interface 93
    input s_axis_bram_93_tlast,
    input s_axis_bram_93_tvalid,
    input [C_INPUT_BRAM_93_DMWIDTH/8-1:0] s_axis_bram_93_tkeep,
    input [C_INPUT_BRAM_93_DMWIDTH/8-1:0] s_axis_bram_93_tstrb,
    input [C_INPUT_BRAM_93_DMWIDTH-1:0] s_axis_bram_93_tdata,
    output s_axis_bram_93_tready,
    input [C_INPUT_BRAM_93_ADDR_WIDTH-1:0] ap_bram_iarg_93_addr0,
    input [C_INPUT_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_din0,
    output [C_INPUT_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_dout0,
    input ap_bram_iarg_93_clk0,
    input ap_bram_iarg_93_rst0,
    input [C_INPUT_BRAM_93_WIDTH/8-1:0] ap_bram_iarg_93_we0,
    input ap_bram_iarg_93_en0,
    input [C_INPUT_BRAM_93_ADDR_WIDTH-1:0] ap_bram_iarg_93_addr1,
    input [C_INPUT_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_din1,
    output [C_INPUT_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_dout1,
    input ap_bram_iarg_93_clk1,
    input ap_bram_iarg_93_rst1,
    input [C_INPUT_BRAM_93_WIDTH/8-1:0] ap_bram_iarg_93_we1,
    input ap_bram_iarg_93_en1,
    //input AXI-Stream to BRAM interface 94
    input s_axis_bram_94_tlast,
    input s_axis_bram_94_tvalid,
    input [C_INPUT_BRAM_94_DMWIDTH/8-1:0] s_axis_bram_94_tkeep,
    input [C_INPUT_BRAM_94_DMWIDTH/8-1:0] s_axis_bram_94_tstrb,
    input [C_INPUT_BRAM_94_DMWIDTH-1:0] s_axis_bram_94_tdata,
    output s_axis_bram_94_tready,
    input [C_INPUT_BRAM_94_ADDR_WIDTH-1:0] ap_bram_iarg_94_addr0,
    input [C_INPUT_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_din0,
    output [C_INPUT_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_dout0,
    input ap_bram_iarg_94_clk0,
    input ap_bram_iarg_94_rst0,
    input [C_INPUT_BRAM_94_WIDTH/8-1:0] ap_bram_iarg_94_we0,
    input ap_bram_iarg_94_en0,
    input [C_INPUT_BRAM_94_ADDR_WIDTH-1:0] ap_bram_iarg_94_addr1,
    input [C_INPUT_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_din1,
    output [C_INPUT_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_dout1,
    input ap_bram_iarg_94_clk1,
    input ap_bram_iarg_94_rst1,
    input [C_INPUT_BRAM_94_WIDTH/8-1:0] ap_bram_iarg_94_we1,
    input ap_bram_iarg_94_en1,
    //input AXI-Stream to BRAM interface 95
    input s_axis_bram_95_tlast,
    input s_axis_bram_95_tvalid,
    input [C_INPUT_BRAM_95_DMWIDTH/8-1:0] s_axis_bram_95_tkeep,
    input [C_INPUT_BRAM_95_DMWIDTH/8-1:0] s_axis_bram_95_tstrb,
    input [C_INPUT_BRAM_95_DMWIDTH-1:0] s_axis_bram_95_tdata,
    output s_axis_bram_95_tready,
    input [C_INPUT_BRAM_95_ADDR_WIDTH-1:0] ap_bram_iarg_95_addr0,
    input [C_INPUT_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_din0,
    output [C_INPUT_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_dout0,
    input ap_bram_iarg_95_clk0,
    input ap_bram_iarg_95_rst0,
    input [C_INPUT_BRAM_95_WIDTH/8-1:0] ap_bram_iarg_95_we0,
    input ap_bram_iarg_95_en0,
    input [C_INPUT_BRAM_95_ADDR_WIDTH-1:0] ap_bram_iarg_95_addr1,
    input [C_INPUT_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_din1,
    output [C_INPUT_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_dout1,
    input ap_bram_iarg_95_clk1,
    input ap_bram_iarg_95_rst1,
    input [C_INPUT_BRAM_95_WIDTH/8-1:0] ap_bram_iarg_95_we1,
    input ap_bram_iarg_95_en1,
    //input AXI-Stream to BRAM interface 96
    input s_axis_bram_96_tlast,
    input s_axis_bram_96_tvalid,
    input [C_INPUT_BRAM_96_DMWIDTH/8-1:0] s_axis_bram_96_tkeep,
    input [C_INPUT_BRAM_96_DMWIDTH/8-1:0] s_axis_bram_96_tstrb,
    input [C_INPUT_BRAM_96_DMWIDTH-1:0] s_axis_bram_96_tdata,
    output s_axis_bram_96_tready,
    input [C_INPUT_BRAM_96_ADDR_WIDTH-1:0] ap_bram_iarg_96_addr0,
    input [C_INPUT_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_din0,
    output [C_INPUT_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_dout0,
    input ap_bram_iarg_96_clk0,
    input ap_bram_iarg_96_rst0,
    input [C_INPUT_BRAM_96_WIDTH/8-1:0] ap_bram_iarg_96_we0,
    input ap_bram_iarg_96_en0,
    input [C_INPUT_BRAM_96_ADDR_WIDTH-1:0] ap_bram_iarg_96_addr1,
    input [C_INPUT_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_din1,
    output [C_INPUT_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_dout1,
    input ap_bram_iarg_96_clk1,
    input ap_bram_iarg_96_rst1,
    input [C_INPUT_BRAM_96_WIDTH/8-1:0] ap_bram_iarg_96_we1,
    input ap_bram_iarg_96_en1,
    //input AXI-Stream to BRAM interface 97
    input s_axis_bram_97_tlast,
    input s_axis_bram_97_tvalid,
    input [C_INPUT_BRAM_97_DMWIDTH/8-1:0] s_axis_bram_97_tkeep,
    input [C_INPUT_BRAM_97_DMWIDTH/8-1:0] s_axis_bram_97_tstrb,
    input [C_INPUT_BRAM_97_DMWIDTH-1:0] s_axis_bram_97_tdata,
    output s_axis_bram_97_tready,
    input [C_INPUT_BRAM_97_ADDR_WIDTH-1:0] ap_bram_iarg_97_addr0,
    input [C_INPUT_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_din0,
    output [C_INPUT_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_dout0,
    input ap_bram_iarg_97_clk0,
    input ap_bram_iarg_97_rst0,
    input [C_INPUT_BRAM_97_WIDTH/8-1:0] ap_bram_iarg_97_we0,
    input ap_bram_iarg_97_en0,
    input [C_INPUT_BRAM_97_ADDR_WIDTH-1:0] ap_bram_iarg_97_addr1,
    input [C_INPUT_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_din1,
    output [C_INPUT_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_dout1,
    input ap_bram_iarg_97_clk1,
    input ap_bram_iarg_97_rst1,
    input [C_INPUT_BRAM_97_WIDTH/8-1:0] ap_bram_iarg_97_we1,
    input ap_bram_iarg_97_en1,
    //input AXI-Stream to BRAM interface 98
    input s_axis_bram_98_tlast,
    input s_axis_bram_98_tvalid,
    input [C_INPUT_BRAM_98_DMWIDTH/8-1:0] s_axis_bram_98_tkeep,
    input [C_INPUT_BRAM_98_DMWIDTH/8-1:0] s_axis_bram_98_tstrb,
    input [C_INPUT_BRAM_98_DMWIDTH-1:0] s_axis_bram_98_tdata,
    output s_axis_bram_98_tready,
    input [C_INPUT_BRAM_98_ADDR_WIDTH-1:0] ap_bram_iarg_98_addr0,
    input [C_INPUT_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_din0,
    output [C_INPUT_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_dout0,
    input ap_bram_iarg_98_clk0,
    input ap_bram_iarg_98_rst0,
    input [C_INPUT_BRAM_98_WIDTH/8-1:0] ap_bram_iarg_98_we0,
    input ap_bram_iarg_98_en0,
    input [C_INPUT_BRAM_98_ADDR_WIDTH-1:0] ap_bram_iarg_98_addr1,
    input [C_INPUT_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_din1,
    output [C_INPUT_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_dout1,
    input ap_bram_iarg_98_clk1,
    input ap_bram_iarg_98_rst1,
    input [C_INPUT_BRAM_98_WIDTH/8-1:0] ap_bram_iarg_98_we1,
    input ap_bram_iarg_98_en1,
    //input AXI-Stream to BRAM interface 99
    input s_axis_bram_99_tlast,
    input s_axis_bram_99_tvalid,
    input [C_INPUT_BRAM_99_DMWIDTH/8-1:0] s_axis_bram_99_tkeep,
    input [C_INPUT_BRAM_99_DMWIDTH/8-1:0] s_axis_bram_99_tstrb,
    input [C_INPUT_BRAM_99_DMWIDTH-1:0] s_axis_bram_99_tdata,
    output s_axis_bram_99_tready,
    input [C_INPUT_BRAM_99_ADDR_WIDTH-1:0] ap_bram_iarg_99_addr0,
    input [C_INPUT_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_din0,
    output [C_INPUT_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_dout0,
    input ap_bram_iarg_99_clk0,
    input ap_bram_iarg_99_rst0,
    input [C_INPUT_BRAM_99_WIDTH/8-1:0] ap_bram_iarg_99_we0,
    input ap_bram_iarg_99_en0,
    input [C_INPUT_BRAM_99_ADDR_WIDTH-1:0] ap_bram_iarg_99_addr1,
    input [C_INPUT_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_din1,
    output [C_INPUT_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_dout1,
    input ap_bram_iarg_99_clk1,
    input ap_bram_iarg_99_rst1,
    input [C_INPUT_BRAM_99_WIDTH/8-1:0] ap_bram_iarg_99_we1,
    input ap_bram_iarg_99_en1,
    //input AXI-Stream to BRAM interface 100
    input s_axis_bram_100_tlast,
    input s_axis_bram_100_tvalid,
    input [C_INPUT_BRAM_100_DMWIDTH/8-1:0] s_axis_bram_100_tkeep,
    input [C_INPUT_BRAM_100_DMWIDTH/8-1:0] s_axis_bram_100_tstrb,
    input [C_INPUT_BRAM_100_DMWIDTH-1:0] s_axis_bram_100_tdata,
    output s_axis_bram_100_tready,
    input [C_INPUT_BRAM_100_ADDR_WIDTH-1:0] ap_bram_iarg_100_addr0,
    input [C_INPUT_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_din0,
    output [C_INPUT_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_dout0,
    input ap_bram_iarg_100_clk0,
    input ap_bram_iarg_100_rst0,
    input [C_INPUT_BRAM_100_WIDTH/8-1:0] ap_bram_iarg_100_we0,
    input ap_bram_iarg_100_en0,
    input [C_INPUT_BRAM_100_ADDR_WIDTH-1:0] ap_bram_iarg_100_addr1,
    input [C_INPUT_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_din1,
    output [C_INPUT_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_dout1,
    input ap_bram_iarg_100_clk1,
    input ap_bram_iarg_100_rst1,
    input [C_INPUT_BRAM_100_WIDTH/8-1:0] ap_bram_iarg_100_we1,
    input ap_bram_iarg_100_en1,
    //input AXI-Stream to BRAM interface 101
    input s_axis_bram_101_tlast,
    input s_axis_bram_101_tvalid,
    input [C_INPUT_BRAM_101_DMWIDTH/8-1:0] s_axis_bram_101_tkeep,
    input [C_INPUT_BRAM_101_DMWIDTH/8-1:0] s_axis_bram_101_tstrb,
    input [C_INPUT_BRAM_101_DMWIDTH-1:0] s_axis_bram_101_tdata,
    output s_axis_bram_101_tready,
    input [C_INPUT_BRAM_101_ADDR_WIDTH-1:0] ap_bram_iarg_101_addr0,
    input [C_INPUT_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_din0,
    output [C_INPUT_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_dout0,
    input ap_bram_iarg_101_clk0,
    input ap_bram_iarg_101_rst0,
    input [C_INPUT_BRAM_101_WIDTH/8-1:0] ap_bram_iarg_101_we0,
    input ap_bram_iarg_101_en0,
    input [C_INPUT_BRAM_101_ADDR_WIDTH-1:0] ap_bram_iarg_101_addr1,
    input [C_INPUT_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_din1,
    output [C_INPUT_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_dout1,
    input ap_bram_iarg_101_clk1,
    input ap_bram_iarg_101_rst1,
    input [C_INPUT_BRAM_101_WIDTH/8-1:0] ap_bram_iarg_101_we1,
    input ap_bram_iarg_101_en1,
    //input AXI-Stream to BRAM interface 102
    input s_axis_bram_102_tlast,
    input s_axis_bram_102_tvalid,
    input [C_INPUT_BRAM_102_DMWIDTH/8-1:0] s_axis_bram_102_tkeep,
    input [C_INPUT_BRAM_102_DMWIDTH/8-1:0] s_axis_bram_102_tstrb,
    input [C_INPUT_BRAM_102_DMWIDTH-1:0] s_axis_bram_102_tdata,
    output s_axis_bram_102_tready,
    input [C_INPUT_BRAM_102_ADDR_WIDTH-1:0] ap_bram_iarg_102_addr0,
    input [C_INPUT_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_din0,
    output [C_INPUT_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_dout0,
    input ap_bram_iarg_102_clk0,
    input ap_bram_iarg_102_rst0,
    input [C_INPUT_BRAM_102_WIDTH/8-1:0] ap_bram_iarg_102_we0,
    input ap_bram_iarg_102_en0,
    input [C_INPUT_BRAM_102_ADDR_WIDTH-1:0] ap_bram_iarg_102_addr1,
    input [C_INPUT_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_din1,
    output [C_INPUT_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_dout1,
    input ap_bram_iarg_102_clk1,
    input ap_bram_iarg_102_rst1,
    input [C_INPUT_BRAM_102_WIDTH/8-1:0] ap_bram_iarg_102_we1,
    input ap_bram_iarg_102_en1,
    //input AXI-Stream to BRAM interface 103
    input s_axis_bram_103_tlast,
    input s_axis_bram_103_tvalid,
    input [C_INPUT_BRAM_103_DMWIDTH/8-1:0] s_axis_bram_103_tkeep,
    input [C_INPUT_BRAM_103_DMWIDTH/8-1:0] s_axis_bram_103_tstrb,
    input [C_INPUT_BRAM_103_DMWIDTH-1:0] s_axis_bram_103_tdata,
    output s_axis_bram_103_tready,
    input [C_INPUT_BRAM_103_ADDR_WIDTH-1:0] ap_bram_iarg_103_addr0,
    input [C_INPUT_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_din0,
    output [C_INPUT_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_dout0,
    input ap_bram_iarg_103_clk0,
    input ap_bram_iarg_103_rst0,
    input [C_INPUT_BRAM_103_WIDTH/8-1:0] ap_bram_iarg_103_we0,
    input ap_bram_iarg_103_en0,
    input [C_INPUT_BRAM_103_ADDR_WIDTH-1:0] ap_bram_iarg_103_addr1,
    input [C_INPUT_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_din1,
    output [C_INPUT_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_dout1,
    input ap_bram_iarg_103_clk1,
    input ap_bram_iarg_103_rst1,
    input [C_INPUT_BRAM_103_WIDTH/8-1:0] ap_bram_iarg_103_we1,
    input ap_bram_iarg_103_en1,
    //input AXI-Stream to BRAM interface 104
    input s_axis_bram_104_tlast,
    input s_axis_bram_104_tvalid,
    input [C_INPUT_BRAM_104_DMWIDTH/8-1:0] s_axis_bram_104_tkeep,
    input [C_INPUT_BRAM_104_DMWIDTH/8-1:0] s_axis_bram_104_tstrb,
    input [C_INPUT_BRAM_104_DMWIDTH-1:0] s_axis_bram_104_tdata,
    output s_axis_bram_104_tready,
    input [C_INPUT_BRAM_104_ADDR_WIDTH-1:0] ap_bram_iarg_104_addr0,
    input [C_INPUT_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_din0,
    output [C_INPUT_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_dout0,
    input ap_bram_iarg_104_clk0,
    input ap_bram_iarg_104_rst0,
    input [C_INPUT_BRAM_104_WIDTH/8-1:0] ap_bram_iarg_104_we0,
    input ap_bram_iarg_104_en0,
    input [C_INPUT_BRAM_104_ADDR_WIDTH-1:0] ap_bram_iarg_104_addr1,
    input [C_INPUT_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_din1,
    output [C_INPUT_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_dout1,
    input ap_bram_iarg_104_clk1,
    input ap_bram_iarg_104_rst1,
    input [C_INPUT_BRAM_104_WIDTH/8-1:0] ap_bram_iarg_104_we1,
    input ap_bram_iarg_104_en1,
    //input AXI-Stream to BRAM interface 105
    input s_axis_bram_105_tlast,
    input s_axis_bram_105_tvalid,
    input [C_INPUT_BRAM_105_DMWIDTH/8-1:0] s_axis_bram_105_tkeep,
    input [C_INPUT_BRAM_105_DMWIDTH/8-1:0] s_axis_bram_105_tstrb,
    input [C_INPUT_BRAM_105_DMWIDTH-1:0] s_axis_bram_105_tdata,
    output s_axis_bram_105_tready,
    input [C_INPUT_BRAM_105_ADDR_WIDTH-1:0] ap_bram_iarg_105_addr0,
    input [C_INPUT_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_din0,
    output [C_INPUT_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_dout0,
    input ap_bram_iarg_105_clk0,
    input ap_bram_iarg_105_rst0,
    input [C_INPUT_BRAM_105_WIDTH/8-1:0] ap_bram_iarg_105_we0,
    input ap_bram_iarg_105_en0,
    input [C_INPUT_BRAM_105_ADDR_WIDTH-1:0] ap_bram_iarg_105_addr1,
    input [C_INPUT_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_din1,
    output [C_INPUT_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_dout1,
    input ap_bram_iarg_105_clk1,
    input ap_bram_iarg_105_rst1,
    input [C_INPUT_BRAM_105_WIDTH/8-1:0] ap_bram_iarg_105_we1,
    input ap_bram_iarg_105_en1,
    //input AXI-Stream to BRAM interface 106
    input s_axis_bram_106_tlast,
    input s_axis_bram_106_tvalid,
    input [C_INPUT_BRAM_106_DMWIDTH/8-1:0] s_axis_bram_106_tkeep,
    input [C_INPUT_BRAM_106_DMWIDTH/8-1:0] s_axis_bram_106_tstrb,
    input [C_INPUT_BRAM_106_DMWIDTH-1:0] s_axis_bram_106_tdata,
    output s_axis_bram_106_tready,
    input [C_INPUT_BRAM_106_ADDR_WIDTH-1:0] ap_bram_iarg_106_addr0,
    input [C_INPUT_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_din0,
    output [C_INPUT_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_dout0,
    input ap_bram_iarg_106_clk0,
    input ap_bram_iarg_106_rst0,
    input [C_INPUT_BRAM_106_WIDTH/8-1:0] ap_bram_iarg_106_we0,
    input ap_bram_iarg_106_en0,
    input [C_INPUT_BRAM_106_ADDR_WIDTH-1:0] ap_bram_iarg_106_addr1,
    input [C_INPUT_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_din1,
    output [C_INPUT_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_dout1,
    input ap_bram_iarg_106_clk1,
    input ap_bram_iarg_106_rst1,
    input [C_INPUT_BRAM_106_WIDTH/8-1:0] ap_bram_iarg_106_we1,
    input ap_bram_iarg_106_en1,
    //input AXI-Stream to BRAM interface 107
    input s_axis_bram_107_tlast,
    input s_axis_bram_107_tvalid,
    input [C_INPUT_BRAM_107_DMWIDTH/8-1:0] s_axis_bram_107_tkeep,
    input [C_INPUT_BRAM_107_DMWIDTH/8-1:0] s_axis_bram_107_tstrb,
    input [C_INPUT_BRAM_107_DMWIDTH-1:0] s_axis_bram_107_tdata,
    output s_axis_bram_107_tready,
    input [C_INPUT_BRAM_107_ADDR_WIDTH-1:0] ap_bram_iarg_107_addr0,
    input [C_INPUT_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_din0,
    output [C_INPUT_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_dout0,
    input ap_bram_iarg_107_clk0,
    input ap_bram_iarg_107_rst0,
    input [C_INPUT_BRAM_107_WIDTH/8-1:0] ap_bram_iarg_107_we0,
    input ap_bram_iarg_107_en0,
    input [C_INPUT_BRAM_107_ADDR_WIDTH-1:0] ap_bram_iarg_107_addr1,
    input [C_INPUT_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_din1,
    output [C_INPUT_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_dout1,
    input ap_bram_iarg_107_clk1,
    input ap_bram_iarg_107_rst1,
    input [C_INPUT_BRAM_107_WIDTH/8-1:0] ap_bram_iarg_107_we1,
    input ap_bram_iarg_107_en1,
    //input AXI-Stream to BRAM interface 108
    input s_axis_bram_108_tlast,
    input s_axis_bram_108_tvalid,
    input [C_INPUT_BRAM_108_DMWIDTH/8-1:0] s_axis_bram_108_tkeep,
    input [C_INPUT_BRAM_108_DMWIDTH/8-1:0] s_axis_bram_108_tstrb,
    input [C_INPUT_BRAM_108_DMWIDTH-1:0] s_axis_bram_108_tdata,
    output s_axis_bram_108_tready,
    input [C_INPUT_BRAM_108_ADDR_WIDTH-1:0] ap_bram_iarg_108_addr0,
    input [C_INPUT_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_din0,
    output [C_INPUT_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_dout0,
    input ap_bram_iarg_108_clk0,
    input ap_bram_iarg_108_rst0,
    input [C_INPUT_BRAM_108_WIDTH/8-1:0] ap_bram_iarg_108_we0,
    input ap_bram_iarg_108_en0,
    input [C_INPUT_BRAM_108_ADDR_WIDTH-1:0] ap_bram_iarg_108_addr1,
    input [C_INPUT_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_din1,
    output [C_INPUT_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_dout1,
    input ap_bram_iarg_108_clk1,
    input ap_bram_iarg_108_rst1,
    input [C_INPUT_BRAM_108_WIDTH/8-1:0] ap_bram_iarg_108_we1,
    input ap_bram_iarg_108_en1,
    //input AXI-Stream to BRAM interface 109
    input s_axis_bram_109_tlast,
    input s_axis_bram_109_tvalid,
    input [C_INPUT_BRAM_109_DMWIDTH/8-1:0] s_axis_bram_109_tkeep,
    input [C_INPUT_BRAM_109_DMWIDTH/8-1:0] s_axis_bram_109_tstrb,
    input [C_INPUT_BRAM_109_DMWIDTH-1:0] s_axis_bram_109_tdata,
    output s_axis_bram_109_tready,
    input [C_INPUT_BRAM_109_ADDR_WIDTH-1:0] ap_bram_iarg_109_addr0,
    input [C_INPUT_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_din0,
    output [C_INPUT_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_dout0,
    input ap_bram_iarg_109_clk0,
    input ap_bram_iarg_109_rst0,
    input [C_INPUT_BRAM_109_WIDTH/8-1:0] ap_bram_iarg_109_we0,
    input ap_bram_iarg_109_en0,
    input [C_INPUT_BRAM_109_ADDR_WIDTH-1:0] ap_bram_iarg_109_addr1,
    input [C_INPUT_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_din1,
    output [C_INPUT_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_dout1,
    input ap_bram_iarg_109_clk1,
    input ap_bram_iarg_109_rst1,
    input [C_INPUT_BRAM_109_WIDTH/8-1:0] ap_bram_iarg_109_we1,
    input ap_bram_iarg_109_en1,
    //input AXI-Stream to BRAM interface 110
    input s_axis_bram_110_tlast,
    input s_axis_bram_110_tvalid,
    input [C_INPUT_BRAM_110_DMWIDTH/8-1:0] s_axis_bram_110_tkeep,
    input [C_INPUT_BRAM_110_DMWIDTH/8-1:0] s_axis_bram_110_tstrb,
    input [C_INPUT_BRAM_110_DMWIDTH-1:0] s_axis_bram_110_tdata,
    output s_axis_bram_110_tready,
    input [C_INPUT_BRAM_110_ADDR_WIDTH-1:0] ap_bram_iarg_110_addr0,
    input [C_INPUT_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_din0,
    output [C_INPUT_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_dout0,
    input ap_bram_iarg_110_clk0,
    input ap_bram_iarg_110_rst0,
    input [C_INPUT_BRAM_110_WIDTH/8-1:0] ap_bram_iarg_110_we0,
    input ap_bram_iarg_110_en0,
    input [C_INPUT_BRAM_110_ADDR_WIDTH-1:0] ap_bram_iarg_110_addr1,
    input [C_INPUT_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_din1,
    output [C_INPUT_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_dout1,
    input ap_bram_iarg_110_clk1,
    input ap_bram_iarg_110_rst1,
    input [C_INPUT_BRAM_110_WIDTH/8-1:0] ap_bram_iarg_110_we1,
    input ap_bram_iarg_110_en1,
    //input AXI-Stream to BRAM interface 111
    input s_axis_bram_111_tlast,
    input s_axis_bram_111_tvalid,
    input [C_INPUT_BRAM_111_DMWIDTH/8-1:0] s_axis_bram_111_tkeep,
    input [C_INPUT_BRAM_111_DMWIDTH/8-1:0] s_axis_bram_111_tstrb,
    input [C_INPUT_BRAM_111_DMWIDTH-1:0] s_axis_bram_111_tdata,
    output s_axis_bram_111_tready,
    input [C_INPUT_BRAM_111_ADDR_WIDTH-1:0] ap_bram_iarg_111_addr0,
    input [C_INPUT_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_din0,
    output [C_INPUT_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_dout0,
    input ap_bram_iarg_111_clk0,
    input ap_bram_iarg_111_rst0,
    input [C_INPUT_BRAM_111_WIDTH/8-1:0] ap_bram_iarg_111_we0,
    input ap_bram_iarg_111_en0,
    input [C_INPUT_BRAM_111_ADDR_WIDTH-1:0] ap_bram_iarg_111_addr1,
    input [C_INPUT_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_din1,
    output [C_INPUT_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_dout1,
    input ap_bram_iarg_111_clk1,
    input ap_bram_iarg_111_rst1,
    input [C_INPUT_BRAM_111_WIDTH/8-1:0] ap_bram_iarg_111_we1,
    input ap_bram_iarg_111_en1,
    //input AXI-Stream to BRAM interface 112
    input s_axis_bram_112_tlast,
    input s_axis_bram_112_tvalid,
    input [C_INPUT_BRAM_112_DMWIDTH/8-1:0] s_axis_bram_112_tkeep,
    input [C_INPUT_BRAM_112_DMWIDTH/8-1:0] s_axis_bram_112_tstrb,
    input [C_INPUT_BRAM_112_DMWIDTH-1:0] s_axis_bram_112_tdata,
    output s_axis_bram_112_tready,
    input [C_INPUT_BRAM_112_ADDR_WIDTH-1:0] ap_bram_iarg_112_addr0,
    input [C_INPUT_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_din0,
    output [C_INPUT_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_dout0,
    input ap_bram_iarg_112_clk0,
    input ap_bram_iarg_112_rst0,
    input [C_INPUT_BRAM_112_WIDTH/8-1:0] ap_bram_iarg_112_we0,
    input ap_bram_iarg_112_en0,
    input [C_INPUT_BRAM_112_ADDR_WIDTH-1:0] ap_bram_iarg_112_addr1,
    input [C_INPUT_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_din1,
    output [C_INPUT_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_dout1,
    input ap_bram_iarg_112_clk1,
    input ap_bram_iarg_112_rst1,
    input [C_INPUT_BRAM_112_WIDTH/8-1:0] ap_bram_iarg_112_we1,
    input ap_bram_iarg_112_en1,
    //input AXI-Stream to BRAM interface 113
    input s_axis_bram_113_tlast,
    input s_axis_bram_113_tvalid,
    input [C_INPUT_BRAM_113_DMWIDTH/8-1:0] s_axis_bram_113_tkeep,
    input [C_INPUT_BRAM_113_DMWIDTH/8-1:0] s_axis_bram_113_tstrb,
    input [C_INPUT_BRAM_113_DMWIDTH-1:0] s_axis_bram_113_tdata,
    output s_axis_bram_113_tready,
    input [C_INPUT_BRAM_113_ADDR_WIDTH-1:0] ap_bram_iarg_113_addr0,
    input [C_INPUT_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_din0,
    output [C_INPUT_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_dout0,
    input ap_bram_iarg_113_clk0,
    input ap_bram_iarg_113_rst0,
    input [C_INPUT_BRAM_113_WIDTH/8-1:0] ap_bram_iarg_113_we0,
    input ap_bram_iarg_113_en0,
    input [C_INPUT_BRAM_113_ADDR_WIDTH-1:0] ap_bram_iarg_113_addr1,
    input [C_INPUT_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_din1,
    output [C_INPUT_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_dout1,
    input ap_bram_iarg_113_clk1,
    input ap_bram_iarg_113_rst1,
    input [C_INPUT_BRAM_113_WIDTH/8-1:0] ap_bram_iarg_113_we1,
    input ap_bram_iarg_113_en1,
    //input AXI-Stream to BRAM interface 114
    input s_axis_bram_114_tlast,
    input s_axis_bram_114_tvalid,
    input [C_INPUT_BRAM_114_DMWIDTH/8-1:0] s_axis_bram_114_tkeep,
    input [C_INPUT_BRAM_114_DMWIDTH/8-1:0] s_axis_bram_114_tstrb,
    input [C_INPUT_BRAM_114_DMWIDTH-1:0] s_axis_bram_114_tdata,
    output s_axis_bram_114_tready,
    input [C_INPUT_BRAM_114_ADDR_WIDTH-1:0] ap_bram_iarg_114_addr0,
    input [C_INPUT_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_din0,
    output [C_INPUT_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_dout0,
    input ap_bram_iarg_114_clk0,
    input ap_bram_iarg_114_rst0,
    input [C_INPUT_BRAM_114_WIDTH/8-1:0] ap_bram_iarg_114_we0,
    input ap_bram_iarg_114_en0,
    input [C_INPUT_BRAM_114_ADDR_WIDTH-1:0] ap_bram_iarg_114_addr1,
    input [C_INPUT_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_din1,
    output [C_INPUT_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_dout1,
    input ap_bram_iarg_114_clk1,
    input ap_bram_iarg_114_rst1,
    input [C_INPUT_BRAM_114_WIDTH/8-1:0] ap_bram_iarg_114_we1,
    input ap_bram_iarg_114_en1,
    //input AXI-Stream to BRAM interface 115
    input s_axis_bram_115_tlast,
    input s_axis_bram_115_tvalid,
    input [C_INPUT_BRAM_115_DMWIDTH/8-1:0] s_axis_bram_115_tkeep,
    input [C_INPUT_BRAM_115_DMWIDTH/8-1:0] s_axis_bram_115_tstrb,
    input [C_INPUT_BRAM_115_DMWIDTH-1:0] s_axis_bram_115_tdata,
    output s_axis_bram_115_tready,
    input [C_INPUT_BRAM_115_ADDR_WIDTH-1:0] ap_bram_iarg_115_addr0,
    input [C_INPUT_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_din0,
    output [C_INPUT_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_dout0,
    input ap_bram_iarg_115_clk0,
    input ap_bram_iarg_115_rst0,
    input [C_INPUT_BRAM_115_WIDTH/8-1:0] ap_bram_iarg_115_we0,
    input ap_bram_iarg_115_en0,
    input [C_INPUT_BRAM_115_ADDR_WIDTH-1:0] ap_bram_iarg_115_addr1,
    input [C_INPUT_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_din1,
    output [C_INPUT_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_dout1,
    input ap_bram_iarg_115_clk1,
    input ap_bram_iarg_115_rst1,
    input [C_INPUT_BRAM_115_WIDTH/8-1:0] ap_bram_iarg_115_we1,
    input ap_bram_iarg_115_en1,
    //input AXI-Stream to BRAM interface 116
    input s_axis_bram_116_tlast,
    input s_axis_bram_116_tvalid,
    input [C_INPUT_BRAM_116_DMWIDTH/8-1:0] s_axis_bram_116_tkeep,
    input [C_INPUT_BRAM_116_DMWIDTH/8-1:0] s_axis_bram_116_tstrb,
    input [C_INPUT_BRAM_116_DMWIDTH-1:0] s_axis_bram_116_tdata,
    output s_axis_bram_116_tready,
    input [C_INPUT_BRAM_116_ADDR_WIDTH-1:0] ap_bram_iarg_116_addr0,
    input [C_INPUT_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_din0,
    output [C_INPUT_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_dout0,
    input ap_bram_iarg_116_clk0,
    input ap_bram_iarg_116_rst0,
    input [C_INPUT_BRAM_116_WIDTH/8-1:0] ap_bram_iarg_116_we0,
    input ap_bram_iarg_116_en0,
    input [C_INPUT_BRAM_116_ADDR_WIDTH-1:0] ap_bram_iarg_116_addr1,
    input [C_INPUT_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_din1,
    output [C_INPUT_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_dout1,
    input ap_bram_iarg_116_clk1,
    input ap_bram_iarg_116_rst1,
    input [C_INPUT_BRAM_116_WIDTH/8-1:0] ap_bram_iarg_116_we1,
    input ap_bram_iarg_116_en1,
    //input AXI-Stream to BRAM interface 117
    input s_axis_bram_117_tlast,
    input s_axis_bram_117_tvalid,
    input [C_INPUT_BRAM_117_DMWIDTH/8-1:0] s_axis_bram_117_tkeep,
    input [C_INPUT_BRAM_117_DMWIDTH/8-1:0] s_axis_bram_117_tstrb,
    input [C_INPUT_BRAM_117_DMWIDTH-1:0] s_axis_bram_117_tdata,
    output s_axis_bram_117_tready,
    input [C_INPUT_BRAM_117_ADDR_WIDTH-1:0] ap_bram_iarg_117_addr0,
    input [C_INPUT_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_din0,
    output [C_INPUT_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_dout0,
    input ap_bram_iarg_117_clk0,
    input ap_bram_iarg_117_rst0,
    input [C_INPUT_BRAM_117_WIDTH/8-1:0] ap_bram_iarg_117_we0,
    input ap_bram_iarg_117_en0,
    input [C_INPUT_BRAM_117_ADDR_WIDTH-1:0] ap_bram_iarg_117_addr1,
    input [C_INPUT_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_din1,
    output [C_INPUT_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_dout1,
    input ap_bram_iarg_117_clk1,
    input ap_bram_iarg_117_rst1,
    input [C_INPUT_BRAM_117_WIDTH/8-1:0] ap_bram_iarg_117_we1,
    input ap_bram_iarg_117_en1,
    //input AXI-Stream to BRAM interface 118
    input s_axis_bram_118_tlast,
    input s_axis_bram_118_tvalid,
    input [C_INPUT_BRAM_118_DMWIDTH/8-1:0] s_axis_bram_118_tkeep,
    input [C_INPUT_BRAM_118_DMWIDTH/8-1:0] s_axis_bram_118_tstrb,
    input [C_INPUT_BRAM_118_DMWIDTH-1:0] s_axis_bram_118_tdata,
    output s_axis_bram_118_tready,
    input [C_INPUT_BRAM_118_ADDR_WIDTH-1:0] ap_bram_iarg_118_addr0,
    input [C_INPUT_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_din0,
    output [C_INPUT_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_dout0,
    input ap_bram_iarg_118_clk0,
    input ap_bram_iarg_118_rst0,
    input [C_INPUT_BRAM_118_WIDTH/8-1:0] ap_bram_iarg_118_we0,
    input ap_bram_iarg_118_en0,
    input [C_INPUT_BRAM_118_ADDR_WIDTH-1:0] ap_bram_iarg_118_addr1,
    input [C_INPUT_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_din1,
    output [C_INPUT_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_dout1,
    input ap_bram_iarg_118_clk1,
    input ap_bram_iarg_118_rst1,
    input [C_INPUT_BRAM_118_WIDTH/8-1:0] ap_bram_iarg_118_we1,
    input ap_bram_iarg_118_en1,
    //input AXI-Stream to BRAM interface 119
    input s_axis_bram_119_tlast,
    input s_axis_bram_119_tvalid,
    input [C_INPUT_BRAM_119_DMWIDTH/8-1:0] s_axis_bram_119_tkeep,
    input [C_INPUT_BRAM_119_DMWIDTH/8-1:0] s_axis_bram_119_tstrb,
    input [C_INPUT_BRAM_119_DMWIDTH-1:0] s_axis_bram_119_tdata,
    output s_axis_bram_119_tready,
    input [C_INPUT_BRAM_119_ADDR_WIDTH-1:0] ap_bram_iarg_119_addr0,
    input [C_INPUT_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_din0,
    output [C_INPUT_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_dout0,
    input ap_bram_iarg_119_clk0,
    input ap_bram_iarg_119_rst0,
    input [C_INPUT_BRAM_119_WIDTH/8-1:0] ap_bram_iarg_119_we0,
    input ap_bram_iarg_119_en0,
    input [C_INPUT_BRAM_119_ADDR_WIDTH-1:0] ap_bram_iarg_119_addr1,
    input [C_INPUT_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_din1,
    output [C_INPUT_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_dout1,
    input ap_bram_iarg_119_clk1,
    input ap_bram_iarg_119_rst1,
    input [C_INPUT_BRAM_119_WIDTH/8-1:0] ap_bram_iarg_119_we1,
    input ap_bram_iarg_119_en1,
    //input AXI-Stream to BRAM interface 120
    input s_axis_bram_120_tlast,
    input s_axis_bram_120_tvalid,
    input [C_INPUT_BRAM_120_DMWIDTH/8-1:0] s_axis_bram_120_tkeep,
    input [C_INPUT_BRAM_120_DMWIDTH/8-1:0] s_axis_bram_120_tstrb,
    input [C_INPUT_BRAM_120_DMWIDTH-1:0] s_axis_bram_120_tdata,
    output s_axis_bram_120_tready,
    input [C_INPUT_BRAM_120_ADDR_WIDTH-1:0] ap_bram_iarg_120_addr0,
    input [C_INPUT_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_din0,
    output [C_INPUT_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_dout0,
    input ap_bram_iarg_120_clk0,
    input ap_bram_iarg_120_rst0,
    input [C_INPUT_BRAM_120_WIDTH/8-1:0] ap_bram_iarg_120_we0,
    input ap_bram_iarg_120_en0,
    input [C_INPUT_BRAM_120_ADDR_WIDTH-1:0] ap_bram_iarg_120_addr1,
    input [C_INPUT_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_din1,
    output [C_INPUT_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_dout1,
    input ap_bram_iarg_120_clk1,
    input ap_bram_iarg_120_rst1,
    input [C_INPUT_BRAM_120_WIDTH/8-1:0] ap_bram_iarg_120_we1,
    input ap_bram_iarg_120_en1,
    //input AXI-Stream to BRAM interface 121
    input s_axis_bram_121_tlast,
    input s_axis_bram_121_tvalid,
    input [C_INPUT_BRAM_121_DMWIDTH/8-1:0] s_axis_bram_121_tkeep,
    input [C_INPUT_BRAM_121_DMWIDTH/8-1:0] s_axis_bram_121_tstrb,
    input [C_INPUT_BRAM_121_DMWIDTH-1:0] s_axis_bram_121_tdata,
    output s_axis_bram_121_tready,
    input [C_INPUT_BRAM_121_ADDR_WIDTH-1:0] ap_bram_iarg_121_addr0,
    input [C_INPUT_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_din0,
    output [C_INPUT_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_dout0,
    input ap_bram_iarg_121_clk0,
    input ap_bram_iarg_121_rst0,
    input [C_INPUT_BRAM_121_WIDTH/8-1:0] ap_bram_iarg_121_we0,
    input ap_bram_iarg_121_en0,
    input [C_INPUT_BRAM_121_ADDR_WIDTH-1:0] ap_bram_iarg_121_addr1,
    input [C_INPUT_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_din1,
    output [C_INPUT_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_dout1,
    input ap_bram_iarg_121_clk1,
    input ap_bram_iarg_121_rst1,
    input [C_INPUT_BRAM_121_WIDTH/8-1:0] ap_bram_iarg_121_we1,
    input ap_bram_iarg_121_en1,
    //input AXI-Stream to BRAM interface 122
    input s_axis_bram_122_tlast,
    input s_axis_bram_122_tvalid,
    input [C_INPUT_BRAM_122_DMWIDTH/8-1:0] s_axis_bram_122_tkeep,
    input [C_INPUT_BRAM_122_DMWIDTH/8-1:0] s_axis_bram_122_tstrb,
    input [C_INPUT_BRAM_122_DMWIDTH-1:0] s_axis_bram_122_tdata,
    output s_axis_bram_122_tready,
    input [C_INPUT_BRAM_122_ADDR_WIDTH-1:0] ap_bram_iarg_122_addr0,
    input [C_INPUT_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_din0,
    output [C_INPUT_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_dout0,
    input ap_bram_iarg_122_clk0,
    input ap_bram_iarg_122_rst0,
    input [C_INPUT_BRAM_122_WIDTH/8-1:0] ap_bram_iarg_122_we0,
    input ap_bram_iarg_122_en0,
    input [C_INPUT_BRAM_122_ADDR_WIDTH-1:0] ap_bram_iarg_122_addr1,
    input [C_INPUT_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_din1,
    output [C_INPUT_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_dout1,
    input ap_bram_iarg_122_clk1,
    input ap_bram_iarg_122_rst1,
    input [C_INPUT_BRAM_122_WIDTH/8-1:0] ap_bram_iarg_122_we1,
    input ap_bram_iarg_122_en1,
    //input AXI-Stream to BRAM interface 123
    input s_axis_bram_123_tlast,
    input s_axis_bram_123_tvalid,
    input [C_INPUT_BRAM_123_DMWIDTH/8-1:0] s_axis_bram_123_tkeep,
    input [C_INPUT_BRAM_123_DMWIDTH/8-1:0] s_axis_bram_123_tstrb,
    input [C_INPUT_BRAM_123_DMWIDTH-1:0] s_axis_bram_123_tdata,
    output s_axis_bram_123_tready,
    input [C_INPUT_BRAM_123_ADDR_WIDTH-1:0] ap_bram_iarg_123_addr0,
    input [C_INPUT_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_din0,
    output [C_INPUT_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_dout0,
    input ap_bram_iarg_123_clk0,
    input ap_bram_iarg_123_rst0,
    input [C_INPUT_BRAM_123_WIDTH/8-1:0] ap_bram_iarg_123_we0,
    input ap_bram_iarg_123_en0,
    input [C_INPUT_BRAM_123_ADDR_WIDTH-1:0] ap_bram_iarg_123_addr1,
    input [C_INPUT_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_din1,
    output [C_INPUT_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_dout1,
    input ap_bram_iarg_123_clk1,
    input ap_bram_iarg_123_rst1,
    input [C_INPUT_BRAM_123_WIDTH/8-1:0] ap_bram_iarg_123_we1,
    input ap_bram_iarg_123_en1,
    //input AXI-Stream to BRAM interface 124
    input s_axis_bram_124_tlast,
    input s_axis_bram_124_tvalid,
    input [C_INPUT_BRAM_124_DMWIDTH/8-1:0] s_axis_bram_124_tkeep,
    input [C_INPUT_BRAM_124_DMWIDTH/8-1:0] s_axis_bram_124_tstrb,
    input [C_INPUT_BRAM_124_DMWIDTH-1:0] s_axis_bram_124_tdata,
    output s_axis_bram_124_tready,
    input [C_INPUT_BRAM_124_ADDR_WIDTH-1:0] ap_bram_iarg_124_addr0,
    input [C_INPUT_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_din0,
    output [C_INPUT_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_dout0,
    input ap_bram_iarg_124_clk0,
    input ap_bram_iarg_124_rst0,
    input [C_INPUT_BRAM_124_WIDTH/8-1:0] ap_bram_iarg_124_we0,
    input ap_bram_iarg_124_en0,
    input [C_INPUT_BRAM_124_ADDR_WIDTH-1:0] ap_bram_iarg_124_addr1,
    input [C_INPUT_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_din1,
    output [C_INPUT_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_dout1,
    input ap_bram_iarg_124_clk1,
    input ap_bram_iarg_124_rst1,
    input [C_INPUT_BRAM_124_WIDTH/8-1:0] ap_bram_iarg_124_we1,
    input ap_bram_iarg_124_en1,
    //input AXI-Stream to BRAM interface 125
    input s_axis_bram_125_tlast,
    input s_axis_bram_125_tvalid,
    input [C_INPUT_BRAM_125_DMWIDTH/8-1:0] s_axis_bram_125_tkeep,
    input [C_INPUT_BRAM_125_DMWIDTH/8-1:0] s_axis_bram_125_tstrb,
    input [C_INPUT_BRAM_125_DMWIDTH-1:0] s_axis_bram_125_tdata,
    output s_axis_bram_125_tready,
    input [C_INPUT_BRAM_125_ADDR_WIDTH-1:0] ap_bram_iarg_125_addr0,
    input [C_INPUT_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_din0,
    output [C_INPUT_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_dout0,
    input ap_bram_iarg_125_clk0,
    input ap_bram_iarg_125_rst0,
    input [C_INPUT_BRAM_125_WIDTH/8-1:0] ap_bram_iarg_125_we0,
    input ap_bram_iarg_125_en0,
    input [C_INPUT_BRAM_125_ADDR_WIDTH-1:0] ap_bram_iarg_125_addr1,
    input [C_INPUT_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_din1,
    output [C_INPUT_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_dout1,
    input ap_bram_iarg_125_clk1,
    input ap_bram_iarg_125_rst1,
    input [C_INPUT_BRAM_125_WIDTH/8-1:0] ap_bram_iarg_125_we1,
    input ap_bram_iarg_125_en1,
    //input AXI-Stream to BRAM interface 126
    input s_axis_bram_126_tlast,
    input s_axis_bram_126_tvalid,
    input [C_INPUT_BRAM_126_DMWIDTH/8-1:0] s_axis_bram_126_tkeep,
    input [C_INPUT_BRAM_126_DMWIDTH/8-1:0] s_axis_bram_126_tstrb,
    input [C_INPUT_BRAM_126_DMWIDTH-1:0] s_axis_bram_126_tdata,
    output s_axis_bram_126_tready,
    input [C_INPUT_BRAM_126_ADDR_WIDTH-1:0] ap_bram_iarg_126_addr0,
    input [C_INPUT_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_din0,
    output [C_INPUT_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_dout0,
    input ap_bram_iarg_126_clk0,
    input ap_bram_iarg_126_rst0,
    input [C_INPUT_BRAM_126_WIDTH/8-1:0] ap_bram_iarg_126_we0,
    input ap_bram_iarg_126_en0,
    input [C_INPUT_BRAM_126_ADDR_WIDTH-1:0] ap_bram_iarg_126_addr1,
    input [C_INPUT_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_din1,
    output [C_INPUT_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_dout1,
    input ap_bram_iarg_126_clk1,
    input ap_bram_iarg_126_rst1,
    input [C_INPUT_BRAM_126_WIDTH/8-1:0] ap_bram_iarg_126_we1,
    input ap_bram_iarg_126_en1,
    //input AXI-Stream to BRAM interface 127
    input s_axis_bram_127_tlast,
    input s_axis_bram_127_tvalid,
    input [C_INPUT_BRAM_127_DMWIDTH/8-1:0] s_axis_bram_127_tkeep,
    input [C_INPUT_BRAM_127_DMWIDTH/8-1:0] s_axis_bram_127_tstrb,
    input [C_INPUT_BRAM_127_DMWIDTH-1:0] s_axis_bram_127_tdata,
    output s_axis_bram_127_tready,
    input [C_INPUT_BRAM_127_ADDR_WIDTH-1:0] ap_bram_iarg_127_addr0,
    input [C_INPUT_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_din0,
    output [C_INPUT_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_dout0,
    input ap_bram_iarg_127_clk0,
    input ap_bram_iarg_127_rst0,
    input [C_INPUT_BRAM_127_WIDTH/8-1:0] ap_bram_iarg_127_we0,
    input ap_bram_iarg_127_en0,
    input [C_INPUT_BRAM_127_ADDR_WIDTH-1:0] ap_bram_iarg_127_addr1,
    input [C_INPUT_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_din1,
    output [C_INPUT_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_dout1,
    input ap_bram_iarg_127_clk1,
    input ap_bram_iarg_127_rst1,
    input [C_INPUT_BRAM_127_WIDTH/8-1:0] ap_bram_iarg_127_we1,
    input ap_bram_iarg_127_en1,
    //-----------------------------------------------------------
    //in-out BRAM AXI-Stream output interface 0
    output m_axis_bramio_0_tlast,
    output m_axis_bramio_0_tvalid,
    output [C_INOUT_BRAM_0_DMWIDTH/8-1:0] m_axis_bramio_0_tkeep,
    output [C_INOUT_BRAM_0_DMWIDTH/8-1:0] m_axis_bramio_0_tstrb,
    output [C_INOUT_BRAM_0_DMWIDTH-1:0] m_axis_bramio_0_tdata,
    input m_axis_bramio_0_tready,
    //in-out BRAM AXI-Stream output interface 1
    output m_axis_bramio_1_tlast,
    output m_axis_bramio_1_tvalid,
    output [C_INOUT_BRAM_1_DMWIDTH/8-1:0] m_axis_bramio_1_tkeep,
    output [C_INOUT_BRAM_1_DMWIDTH/8-1:0] m_axis_bramio_1_tstrb,
    output [C_INOUT_BRAM_1_DMWIDTH-1:0] m_axis_bramio_1_tdata,
    input m_axis_bramio_1_tready,
    //in-out BRAM AXI-Stream output interface 2
    output m_axis_bramio_2_tlast,
    output m_axis_bramio_2_tvalid,
    output [C_INOUT_BRAM_2_DMWIDTH/8-1:0] m_axis_bramio_2_tkeep,
    output [C_INOUT_BRAM_2_DMWIDTH/8-1:0] m_axis_bramio_2_tstrb,
    output [C_INOUT_BRAM_2_DMWIDTH-1:0] m_axis_bramio_2_tdata,
    input m_axis_bramio_2_tready,
    //in-out BRAM AXI-Stream output interface 3
    output m_axis_bramio_3_tlast,
    output m_axis_bramio_3_tvalid,
    output [C_INOUT_BRAM_3_DMWIDTH/8-1:0] m_axis_bramio_3_tkeep,
    output [C_INOUT_BRAM_3_DMWIDTH/8-1:0] m_axis_bramio_3_tstrb,
    output [C_INOUT_BRAM_3_DMWIDTH-1:0] m_axis_bramio_3_tdata,
    input m_axis_bramio_3_tready,
    //in-out BRAM AXI-Stream output interface 4
    output m_axis_bramio_4_tlast,
    output m_axis_bramio_4_tvalid,
    output [C_INOUT_BRAM_4_DMWIDTH/8-1:0] m_axis_bramio_4_tkeep,
    output [C_INOUT_BRAM_4_DMWIDTH/8-1:0] m_axis_bramio_4_tstrb,
    output [C_INOUT_BRAM_4_DMWIDTH-1:0] m_axis_bramio_4_tdata,
    input m_axis_bramio_4_tready,
    //in-out BRAM AXI-Stream output interface 5
    output m_axis_bramio_5_tlast,
    output m_axis_bramio_5_tvalid,
    output [C_INOUT_BRAM_5_DMWIDTH/8-1:0] m_axis_bramio_5_tkeep,
    output [C_INOUT_BRAM_5_DMWIDTH/8-1:0] m_axis_bramio_5_tstrb,
    output [C_INOUT_BRAM_5_DMWIDTH-1:0] m_axis_bramio_5_tdata,
    input m_axis_bramio_5_tready,
    //in-out BRAM AXI-Stream output interface 6
    output m_axis_bramio_6_tlast,
    output m_axis_bramio_6_tvalid,
    output [C_INOUT_BRAM_6_DMWIDTH/8-1:0] m_axis_bramio_6_tkeep,
    output [C_INOUT_BRAM_6_DMWIDTH/8-1:0] m_axis_bramio_6_tstrb,
    output [C_INOUT_BRAM_6_DMWIDTH-1:0] m_axis_bramio_6_tdata,
    input m_axis_bramio_6_tready,
    //in-out BRAM AXI-Stream output interface 7
    output m_axis_bramio_7_tlast,
    output m_axis_bramio_7_tvalid,
    output [C_INOUT_BRAM_7_DMWIDTH/8-1:0] m_axis_bramio_7_tkeep,
    output [C_INOUT_BRAM_7_DMWIDTH/8-1:0] m_axis_bramio_7_tstrb,
    output [C_INOUT_BRAM_7_DMWIDTH-1:0] m_axis_bramio_7_tdata,
    input m_axis_bramio_7_tready,
    //in-out BRAM AXI-Stream output interface 8
    output m_axis_bramio_8_tlast,
    output m_axis_bramio_8_tvalid,
    output [C_INOUT_BRAM_8_DMWIDTH/8-1:0] m_axis_bramio_8_tkeep,
    output [C_INOUT_BRAM_8_DMWIDTH/8-1:0] m_axis_bramio_8_tstrb,
    output [C_INOUT_BRAM_8_DMWIDTH-1:0] m_axis_bramio_8_tdata,
    input m_axis_bramio_8_tready,
    //in-out BRAM AXI-Stream output interface 9
    output m_axis_bramio_9_tlast,
    output m_axis_bramio_9_tvalid,
    output [C_INOUT_BRAM_9_DMWIDTH/8-1:0] m_axis_bramio_9_tkeep,
    output [C_INOUT_BRAM_9_DMWIDTH/8-1:0] m_axis_bramio_9_tstrb,
    output [C_INOUT_BRAM_9_DMWIDTH-1:0] m_axis_bramio_9_tdata,
    input m_axis_bramio_9_tready,
    //in-out BRAM AXI-Stream output interface 10
    output m_axis_bramio_10_tlast,
    output m_axis_bramio_10_tvalid,
    output [C_INOUT_BRAM_10_DMWIDTH/8-1:0] m_axis_bramio_10_tkeep,
    output [C_INOUT_BRAM_10_DMWIDTH/8-1:0] m_axis_bramio_10_tstrb,
    output [C_INOUT_BRAM_10_DMWIDTH-1:0] m_axis_bramio_10_tdata,
    input m_axis_bramio_10_tready,
    //in-out BRAM AXI-Stream output interface 11
    output m_axis_bramio_11_tlast,
    output m_axis_bramio_11_tvalid,
    output [C_INOUT_BRAM_11_DMWIDTH/8-1:0] m_axis_bramio_11_tkeep,
    output [C_INOUT_BRAM_11_DMWIDTH/8-1:0] m_axis_bramio_11_tstrb,
    output [C_INOUT_BRAM_11_DMWIDTH-1:0] m_axis_bramio_11_tdata,
    input m_axis_bramio_11_tready,
    //in-out BRAM AXI-Stream output interface 12
    output m_axis_bramio_12_tlast,
    output m_axis_bramio_12_tvalid,
    output [C_INOUT_BRAM_12_DMWIDTH/8-1:0] m_axis_bramio_12_tkeep,
    output [C_INOUT_BRAM_12_DMWIDTH/8-1:0] m_axis_bramio_12_tstrb,
    output [C_INOUT_BRAM_12_DMWIDTH-1:0] m_axis_bramio_12_tdata,
    input m_axis_bramio_12_tready,
    //in-out BRAM AXI-Stream output interface 13
    output m_axis_bramio_13_tlast,
    output m_axis_bramio_13_tvalid,
    output [C_INOUT_BRAM_13_DMWIDTH/8-1:0] m_axis_bramio_13_tkeep,
    output [C_INOUT_BRAM_13_DMWIDTH/8-1:0] m_axis_bramio_13_tstrb,
    output [C_INOUT_BRAM_13_DMWIDTH-1:0] m_axis_bramio_13_tdata,
    input m_axis_bramio_13_tready,
    //in-out BRAM AXI-Stream output interface 14
    output m_axis_bramio_14_tlast,
    output m_axis_bramio_14_tvalid,
    output [C_INOUT_BRAM_14_DMWIDTH/8-1:0] m_axis_bramio_14_tkeep,
    output [C_INOUT_BRAM_14_DMWIDTH/8-1:0] m_axis_bramio_14_tstrb,
    output [C_INOUT_BRAM_14_DMWIDTH-1:0] m_axis_bramio_14_tdata,
    input m_axis_bramio_14_tready,
    //in-out BRAM AXI-Stream output interface 15
    output m_axis_bramio_15_tlast,
    output m_axis_bramio_15_tvalid,
    output [C_INOUT_BRAM_15_DMWIDTH/8-1:0] m_axis_bramio_15_tkeep,
    output [C_INOUT_BRAM_15_DMWIDTH/8-1:0] m_axis_bramio_15_tstrb,
    output [C_INOUT_BRAM_15_DMWIDTH-1:0] m_axis_bramio_15_tdata,
    input m_axis_bramio_15_tready,
    //in-out BRAM AXI-Stream output interface 16
    output m_axis_bramio_16_tlast,
    output m_axis_bramio_16_tvalid,
    output [C_INOUT_BRAM_16_DMWIDTH/8-1:0] m_axis_bramio_16_tkeep,
    output [C_INOUT_BRAM_16_DMWIDTH/8-1:0] m_axis_bramio_16_tstrb,
    output [C_INOUT_BRAM_16_DMWIDTH-1:0] m_axis_bramio_16_tdata,
    input m_axis_bramio_16_tready,
    //in-out BRAM AXI-Stream output interface 17
    output m_axis_bramio_17_tlast,
    output m_axis_bramio_17_tvalid,
    output [C_INOUT_BRAM_17_DMWIDTH/8-1:0] m_axis_bramio_17_tkeep,
    output [C_INOUT_BRAM_17_DMWIDTH/8-1:0] m_axis_bramio_17_tstrb,
    output [C_INOUT_BRAM_17_DMWIDTH-1:0] m_axis_bramio_17_tdata,
    input m_axis_bramio_17_tready,
    //in-out BRAM AXI-Stream output interface 18
    output m_axis_bramio_18_tlast,
    output m_axis_bramio_18_tvalid,
    output [C_INOUT_BRAM_18_DMWIDTH/8-1:0] m_axis_bramio_18_tkeep,
    output [C_INOUT_BRAM_18_DMWIDTH/8-1:0] m_axis_bramio_18_tstrb,
    output [C_INOUT_BRAM_18_DMWIDTH-1:0] m_axis_bramio_18_tdata,
    input m_axis_bramio_18_tready,
    //in-out BRAM AXI-Stream output interface 19
    output m_axis_bramio_19_tlast,
    output m_axis_bramio_19_tvalid,
    output [C_INOUT_BRAM_19_DMWIDTH/8-1:0] m_axis_bramio_19_tkeep,
    output [C_INOUT_BRAM_19_DMWIDTH/8-1:0] m_axis_bramio_19_tstrb,
    output [C_INOUT_BRAM_19_DMWIDTH-1:0] m_axis_bramio_19_tdata,
    input m_axis_bramio_19_tready,
    //in-out BRAM AXI-Stream output interface 20
    output m_axis_bramio_20_tlast,
    output m_axis_bramio_20_tvalid,
    output [C_INOUT_BRAM_20_DMWIDTH/8-1:0] m_axis_bramio_20_tkeep,
    output [C_INOUT_BRAM_20_DMWIDTH/8-1:0] m_axis_bramio_20_tstrb,
    output [C_INOUT_BRAM_20_DMWIDTH-1:0] m_axis_bramio_20_tdata,
    input m_axis_bramio_20_tready,
    //in-out BRAM AXI-Stream output interface 21
    output m_axis_bramio_21_tlast,
    output m_axis_bramio_21_tvalid,
    output [C_INOUT_BRAM_21_DMWIDTH/8-1:0] m_axis_bramio_21_tkeep,
    output [C_INOUT_BRAM_21_DMWIDTH/8-1:0] m_axis_bramio_21_tstrb,
    output [C_INOUT_BRAM_21_DMWIDTH-1:0] m_axis_bramio_21_tdata,
    input m_axis_bramio_21_tready,
    //in-out BRAM AXI-Stream output interface 22
    output m_axis_bramio_22_tlast,
    output m_axis_bramio_22_tvalid,
    output [C_INOUT_BRAM_22_DMWIDTH/8-1:0] m_axis_bramio_22_tkeep,
    output [C_INOUT_BRAM_22_DMWIDTH/8-1:0] m_axis_bramio_22_tstrb,
    output [C_INOUT_BRAM_22_DMWIDTH-1:0] m_axis_bramio_22_tdata,
    input m_axis_bramio_22_tready,
    //in-out BRAM AXI-Stream output interface 23
    output m_axis_bramio_23_tlast,
    output m_axis_bramio_23_tvalid,
    output [C_INOUT_BRAM_23_DMWIDTH/8-1:0] m_axis_bramio_23_tkeep,
    output [C_INOUT_BRAM_23_DMWIDTH/8-1:0] m_axis_bramio_23_tstrb,
    output [C_INOUT_BRAM_23_DMWIDTH-1:0] m_axis_bramio_23_tdata,
    input m_axis_bramio_23_tready,
    //in-out BRAM AXI-Stream output interface 24
    output m_axis_bramio_24_tlast,
    output m_axis_bramio_24_tvalid,
    output [C_INOUT_BRAM_24_DMWIDTH/8-1:0] m_axis_bramio_24_tkeep,
    output [C_INOUT_BRAM_24_DMWIDTH/8-1:0] m_axis_bramio_24_tstrb,
    output [C_INOUT_BRAM_24_DMWIDTH-1:0] m_axis_bramio_24_tdata,
    input m_axis_bramio_24_tready,
    //in-out BRAM AXI-Stream output interface 25
    output m_axis_bramio_25_tlast,
    output m_axis_bramio_25_tvalid,
    output [C_INOUT_BRAM_25_DMWIDTH/8-1:0] m_axis_bramio_25_tkeep,
    output [C_INOUT_BRAM_25_DMWIDTH/8-1:0] m_axis_bramio_25_tstrb,
    output [C_INOUT_BRAM_25_DMWIDTH-1:0] m_axis_bramio_25_tdata,
    input m_axis_bramio_25_tready,
    //in-out BRAM AXI-Stream output interface 26
    output m_axis_bramio_26_tlast,
    output m_axis_bramio_26_tvalid,
    output [C_INOUT_BRAM_26_DMWIDTH/8-1:0] m_axis_bramio_26_tkeep,
    output [C_INOUT_BRAM_26_DMWIDTH/8-1:0] m_axis_bramio_26_tstrb,
    output [C_INOUT_BRAM_26_DMWIDTH-1:0] m_axis_bramio_26_tdata,
    input m_axis_bramio_26_tready,
    //in-out BRAM AXI-Stream output interface 27
    output m_axis_bramio_27_tlast,
    output m_axis_bramio_27_tvalid,
    output [C_INOUT_BRAM_27_DMWIDTH/8-1:0] m_axis_bramio_27_tkeep,
    output [C_INOUT_BRAM_27_DMWIDTH/8-1:0] m_axis_bramio_27_tstrb,
    output [C_INOUT_BRAM_27_DMWIDTH-1:0] m_axis_bramio_27_tdata,
    input m_axis_bramio_27_tready,
    //in-out BRAM AXI-Stream output interface 28
    output m_axis_bramio_28_tlast,
    output m_axis_bramio_28_tvalid,
    output [C_INOUT_BRAM_28_DMWIDTH/8-1:0] m_axis_bramio_28_tkeep,
    output [C_INOUT_BRAM_28_DMWIDTH/8-1:0] m_axis_bramio_28_tstrb,
    output [C_INOUT_BRAM_28_DMWIDTH-1:0] m_axis_bramio_28_tdata,
    input m_axis_bramio_28_tready,
    //in-out BRAM AXI-Stream output interface 29
    output m_axis_bramio_29_tlast,
    output m_axis_bramio_29_tvalid,
    output [C_INOUT_BRAM_29_DMWIDTH/8-1:0] m_axis_bramio_29_tkeep,
    output [C_INOUT_BRAM_29_DMWIDTH/8-1:0] m_axis_bramio_29_tstrb,
    output [C_INOUT_BRAM_29_DMWIDTH-1:0] m_axis_bramio_29_tdata,
    input m_axis_bramio_29_tready,
    //in-out BRAM AXI-Stream output interface 30
    output m_axis_bramio_30_tlast,
    output m_axis_bramio_30_tvalid,
    output [C_INOUT_BRAM_30_DMWIDTH/8-1:0] m_axis_bramio_30_tkeep,
    output [C_INOUT_BRAM_30_DMWIDTH/8-1:0] m_axis_bramio_30_tstrb,
    output [C_INOUT_BRAM_30_DMWIDTH-1:0] m_axis_bramio_30_tdata,
    input m_axis_bramio_30_tready,
    //in-out BRAM AXI-Stream output interface 31
    output m_axis_bramio_31_tlast,
    output m_axis_bramio_31_tvalid,
    output [C_INOUT_BRAM_31_DMWIDTH/8-1:0] m_axis_bramio_31_tkeep,
    output [C_INOUT_BRAM_31_DMWIDTH/8-1:0] m_axis_bramio_31_tstrb,
    output [C_INOUT_BRAM_31_DMWIDTH-1:0] m_axis_bramio_31_tdata,
    input m_axis_bramio_31_tready,
    //in-out BRAM AXI-Stream output interface 32
    output m_axis_bramio_32_tlast,
    output m_axis_bramio_32_tvalid,
    output [C_INOUT_BRAM_32_DMWIDTH/8-1:0] m_axis_bramio_32_tkeep,
    output [C_INOUT_BRAM_32_DMWIDTH/8-1:0] m_axis_bramio_32_tstrb,
    output [C_INOUT_BRAM_32_DMWIDTH-1:0] m_axis_bramio_32_tdata,
    input m_axis_bramio_32_tready,
    //in-out BRAM AXI-Stream output interface 33
    output m_axis_bramio_33_tlast,
    output m_axis_bramio_33_tvalid,
    output [C_INOUT_BRAM_33_DMWIDTH/8-1:0] m_axis_bramio_33_tkeep,
    output [C_INOUT_BRAM_33_DMWIDTH/8-1:0] m_axis_bramio_33_tstrb,
    output [C_INOUT_BRAM_33_DMWIDTH-1:0] m_axis_bramio_33_tdata,
    input m_axis_bramio_33_tready,
    //in-out BRAM AXI-Stream output interface 34
    output m_axis_bramio_34_tlast,
    output m_axis_bramio_34_tvalid,
    output [C_INOUT_BRAM_34_DMWIDTH/8-1:0] m_axis_bramio_34_tkeep,
    output [C_INOUT_BRAM_34_DMWIDTH/8-1:0] m_axis_bramio_34_tstrb,
    output [C_INOUT_BRAM_34_DMWIDTH-1:0] m_axis_bramio_34_tdata,
    input m_axis_bramio_34_tready,
    //in-out BRAM AXI-Stream output interface 35
    output m_axis_bramio_35_tlast,
    output m_axis_bramio_35_tvalid,
    output [C_INOUT_BRAM_35_DMWIDTH/8-1:0] m_axis_bramio_35_tkeep,
    output [C_INOUT_BRAM_35_DMWIDTH/8-1:0] m_axis_bramio_35_tstrb,
    output [C_INOUT_BRAM_35_DMWIDTH-1:0] m_axis_bramio_35_tdata,
    input m_axis_bramio_35_tready,
    //in-out BRAM AXI-Stream output interface 36
    output m_axis_bramio_36_tlast,
    output m_axis_bramio_36_tvalid,
    output [C_INOUT_BRAM_36_DMWIDTH/8-1:0] m_axis_bramio_36_tkeep,
    output [C_INOUT_BRAM_36_DMWIDTH/8-1:0] m_axis_bramio_36_tstrb,
    output [C_INOUT_BRAM_36_DMWIDTH-1:0] m_axis_bramio_36_tdata,
    input m_axis_bramio_36_tready,
    //in-out BRAM AXI-Stream output interface 37
    output m_axis_bramio_37_tlast,
    output m_axis_bramio_37_tvalid,
    output [C_INOUT_BRAM_37_DMWIDTH/8-1:0] m_axis_bramio_37_tkeep,
    output [C_INOUT_BRAM_37_DMWIDTH/8-1:0] m_axis_bramio_37_tstrb,
    output [C_INOUT_BRAM_37_DMWIDTH-1:0] m_axis_bramio_37_tdata,
    input m_axis_bramio_37_tready,
    //in-out BRAM AXI-Stream output interface 38
    output m_axis_bramio_38_tlast,
    output m_axis_bramio_38_tvalid,
    output [C_INOUT_BRAM_38_DMWIDTH/8-1:0] m_axis_bramio_38_tkeep,
    output [C_INOUT_BRAM_38_DMWIDTH/8-1:0] m_axis_bramio_38_tstrb,
    output [C_INOUT_BRAM_38_DMWIDTH-1:0] m_axis_bramio_38_tdata,
    input m_axis_bramio_38_tready,
    //in-out BRAM AXI-Stream output interface 39
    output m_axis_bramio_39_tlast,
    output m_axis_bramio_39_tvalid,
    output [C_INOUT_BRAM_39_DMWIDTH/8-1:0] m_axis_bramio_39_tkeep,
    output [C_INOUT_BRAM_39_DMWIDTH/8-1:0] m_axis_bramio_39_tstrb,
    output [C_INOUT_BRAM_39_DMWIDTH-1:0] m_axis_bramio_39_tdata,
    input m_axis_bramio_39_tready,
    //in-out BRAM AXI-Stream output interface 40
    output m_axis_bramio_40_tlast,
    output m_axis_bramio_40_tvalid,
    output [C_INOUT_BRAM_40_DMWIDTH/8-1:0] m_axis_bramio_40_tkeep,
    output [C_INOUT_BRAM_40_DMWIDTH/8-1:0] m_axis_bramio_40_tstrb,
    output [C_INOUT_BRAM_40_DMWIDTH-1:0] m_axis_bramio_40_tdata,
    input m_axis_bramio_40_tready,
    //in-out BRAM AXI-Stream output interface 41
    output m_axis_bramio_41_tlast,
    output m_axis_bramio_41_tvalid,
    output [C_INOUT_BRAM_41_DMWIDTH/8-1:0] m_axis_bramio_41_tkeep,
    output [C_INOUT_BRAM_41_DMWIDTH/8-1:0] m_axis_bramio_41_tstrb,
    output [C_INOUT_BRAM_41_DMWIDTH-1:0] m_axis_bramio_41_tdata,
    input m_axis_bramio_41_tready,
    //in-out BRAM AXI-Stream output interface 42
    output m_axis_bramio_42_tlast,
    output m_axis_bramio_42_tvalid,
    output [C_INOUT_BRAM_42_DMWIDTH/8-1:0] m_axis_bramio_42_tkeep,
    output [C_INOUT_BRAM_42_DMWIDTH/8-1:0] m_axis_bramio_42_tstrb,
    output [C_INOUT_BRAM_42_DMWIDTH-1:0] m_axis_bramio_42_tdata,
    input m_axis_bramio_42_tready,
    //in-out BRAM AXI-Stream output interface 43
    output m_axis_bramio_43_tlast,
    output m_axis_bramio_43_tvalid,
    output [C_INOUT_BRAM_43_DMWIDTH/8-1:0] m_axis_bramio_43_tkeep,
    output [C_INOUT_BRAM_43_DMWIDTH/8-1:0] m_axis_bramio_43_tstrb,
    output [C_INOUT_BRAM_43_DMWIDTH-1:0] m_axis_bramio_43_tdata,
    input m_axis_bramio_43_tready,
    //in-out BRAM AXI-Stream output interface 44
    output m_axis_bramio_44_tlast,
    output m_axis_bramio_44_tvalid,
    output [C_INOUT_BRAM_44_DMWIDTH/8-1:0] m_axis_bramio_44_tkeep,
    output [C_INOUT_BRAM_44_DMWIDTH/8-1:0] m_axis_bramio_44_tstrb,
    output [C_INOUT_BRAM_44_DMWIDTH-1:0] m_axis_bramio_44_tdata,
    input m_axis_bramio_44_tready,
    //in-out BRAM AXI-Stream output interface 45
    output m_axis_bramio_45_tlast,
    output m_axis_bramio_45_tvalid,
    output [C_INOUT_BRAM_45_DMWIDTH/8-1:0] m_axis_bramio_45_tkeep,
    output [C_INOUT_BRAM_45_DMWIDTH/8-1:0] m_axis_bramio_45_tstrb,
    output [C_INOUT_BRAM_45_DMWIDTH-1:0] m_axis_bramio_45_tdata,
    input m_axis_bramio_45_tready,
    //in-out BRAM AXI-Stream output interface 46
    output m_axis_bramio_46_tlast,
    output m_axis_bramio_46_tvalid,
    output [C_INOUT_BRAM_46_DMWIDTH/8-1:0] m_axis_bramio_46_tkeep,
    output [C_INOUT_BRAM_46_DMWIDTH/8-1:0] m_axis_bramio_46_tstrb,
    output [C_INOUT_BRAM_46_DMWIDTH-1:0] m_axis_bramio_46_tdata,
    input m_axis_bramio_46_tready,
    //in-out BRAM AXI-Stream output interface 47
    output m_axis_bramio_47_tlast,
    output m_axis_bramio_47_tvalid,
    output [C_INOUT_BRAM_47_DMWIDTH/8-1:0] m_axis_bramio_47_tkeep,
    output [C_INOUT_BRAM_47_DMWIDTH/8-1:0] m_axis_bramio_47_tstrb,
    output [C_INOUT_BRAM_47_DMWIDTH-1:0] m_axis_bramio_47_tdata,
    input m_axis_bramio_47_tready,
    //in-out BRAM AXI-Stream output interface 48
    output m_axis_bramio_48_tlast,
    output m_axis_bramio_48_tvalid,
    output [C_INOUT_BRAM_48_DMWIDTH/8-1:0] m_axis_bramio_48_tkeep,
    output [C_INOUT_BRAM_48_DMWIDTH/8-1:0] m_axis_bramio_48_tstrb,
    output [C_INOUT_BRAM_48_DMWIDTH-1:0] m_axis_bramio_48_tdata,
    input m_axis_bramio_48_tready,
    //in-out BRAM AXI-Stream output interface 49
    output m_axis_bramio_49_tlast,
    output m_axis_bramio_49_tvalid,
    output [C_INOUT_BRAM_49_DMWIDTH/8-1:0] m_axis_bramio_49_tkeep,
    output [C_INOUT_BRAM_49_DMWIDTH/8-1:0] m_axis_bramio_49_tstrb,
    output [C_INOUT_BRAM_49_DMWIDTH-1:0] m_axis_bramio_49_tdata,
    input m_axis_bramio_49_tready,
    //in-out BRAM AXI-Stream output interface 50
    output m_axis_bramio_50_tlast,
    output m_axis_bramio_50_tvalid,
    output [C_INOUT_BRAM_50_DMWIDTH/8-1:0] m_axis_bramio_50_tkeep,
    output [C_INOUT_BRAM_50_DMWIDTH/8-1:0] m_axis_bramio_50_tstrb,
    output [C_INOUT_BRAM_50_DMWIDTH-1:0] m_axis_bramio_50_tdata,
    input m_axis_bramio_50_tready,
    //in-out BRAM AXI-Stream output interface 51
    output m_axis_bramio_51_tlast,
    output m_axis_bramio_51_tvalid,
    output [C_INOUT_BRAM_51_DMWIDTH/8-1:0] m_axis_bramio_51_tkeep,
    output [C_INOUT_BRAM_51_DMWIDTH/8-1:0] m_axis_bramio_51_tstrb,
    output [C_INOUT_BRAM_51_DMWIDTH-1:0] m_axis_bramio_51_tdata,
    input m_axis_bramio_51_tready,
    //in-out BRAM AXI-Stream output interface 52
    output m_axis_bramio_52_tlast,
    output m_axis_bramio_52_tvalid,
    output [C_INOUT_BRAM_52_DMWIDTH/8-1:0] m_axis_bramio_52_tkeep,
    output [C_INOUT_BRAM_52_DMWIDTH/8-1:0] m_axis_bramio_52_tstrb,
    output [C_INOUT_BRAM_52_DMWIDTH-1:0] m_axis_bramio_52_tdata,
    input m_axis_bramio_52_tready,
    //in-out BRAM AXI-Stream output interface 53
    output m_axis_bramio_53_tlast,
    output m_axis_bramio_53_tvalid,
    output [C_INOUT_BRAM_53_DMWIDTH/8-1:0] m_axis_bramio_53_tkeep,
    output [C_INOUT_BRAM_53_DMWIDTH/8-1:0] m_axis_bramio_53_tstrb,
    output [C_INOUT_BRAM_53_DMWIDTH-1:0] m_axis_bramio_53_tdata,
    input m_axis_bramio_53_tready,
    //in-out BRAM AXI-Stream output interface 54
    output m_axis_bramio_54_tlast,
    output m_axis_bramio_54_tvalid,
    output [C_INOUT_BRAM_54_DMWIDTH/8-1:0] m_axis_bramio_54_tkeep,
    output [C_INOUT_BRAM_54_DMWIDTH/8-1:0] m_axis_bramio_54_tstrb,
    output [C_INOUT_BRAM_54_DMWIDTH-1:0] m_axis_bramio_54_tdata,
    input m_axis_bramio_54_tready,
    //in-out BRAM AXI-Stream output interface 55
    output m_axis_bramio_55_tlast,
    output m_axis_bramio_55_tvalid,
    output [C_INOUT_BRAM_55_DMWIDTH/8-1:0] m_axis_bramio_55_tkeep,
    output [C_INOUT_BRAM_55_DMWIDTH/8-1:0] m_axis_bramio_55_tstrb,
    output [C_INOUT_BRAM_55_DMWIDTH-1:0] m_axis_bramio_55_tdata,
    input m_axis_bramio_55_tready,
    //in-out BRAM AXI-Stream output interface 56
    output m_axis_bramio_56_tlast,
    output m_axis_bramio_56_tvalid,
    output [C_INOUT_BRAM_56_DMWIDTH/8-1:0] m_axis_bramio_56_tkeep,
    output [C_INOUT_BRAM_56_DMWIDTH/8-1:0] m_axis_bramio_56_tstrb,
    output [C_INOUT_BRAM_56_DMWIDTH-1:0] m_axis_bramio_56_tdata,
    input m_axis_bramio_56_tready,
    //in-out BRAM AXI-Stream output interface 57
    output m_axis_bramio_57_tlast,
    output m_axis_bramio_57_tvalid,
    output [C_INOUT_BRAM_57_DMWIDTH/8-1:0] m_axis_bramio_57_tkeep,
    output [C_INOUT_BRAM_57_DMWIDTH/8-1:0] m_axis_bramio_57_tstrb,
    output [C_INOUT_BRAM_57_DMWIDTH-1:0] m_axis_bramio_57_tdata,
    input m_axis_bramio_57_tready,
    //in-out BRAM AXI-Stream output interface 58
    output m_axis_bramio_58_tlast,
    output m_axis_bramio_58_tvalid,
    output [C_INOUT_BRAM_58_DMWIDTH/8-1:0] m_axis_bramio_58_tkeep,
    output [C_INOUT_BRAM_58_DMWIDTH/8-1:0] m_axis_bramio_58_tstrb,
    output [C_INOUT_BRAM_58_DMWIDTH-1:0] m_axis_bramio_58_tdata,
    input m_axis_bramio_58_tready,
    //in-out BRAM AXI-Stream output interface 59
    output m_axis_bramio_59_tlast,
    output m_axis_bramio_59_tvalid,
    output [C_INOUT_BRAM_59_DMWIDTH/8-1:0] m_axis_bramio_59_tkeep,
    output [C_INOUT_BRAM_59_DMWIDTH/8-1:0] m_axis_bramio_59_tstrb,
    output [C_INOUT_BRAM_59_DMWIDTH-1:0] m_axis_bramio_59_tdata,
    input m_axis_bramio_59_tready,
    //in-out BRAM AXI-Stream output interface 60
    output m_axis_bramio_60_tlast,
    output m_axis_bramio_60_tvalid,
    output [C_INOUT_BRAM_60_DMWIDTH/8-1:0] m_axis_bramio_60_tkeep,
    output [C_INOUT_BRAM_60_DMWIDTH/8-1:0] m_axis_bramio_60_tstrb,
    output [C_INOUT_BRAM_60_DMWIDTH-1:0] m_axis_bramio_60_tdata,
    input m_axis_bramio_60_tready,
    //in-out BRAM AXI-Stream output interface 61
    output m_axis_bramio_61_tlast,
    output m_axis_bramio_61_tvalid,
    output [C_INOUT_BRAM_61_DMWIDTH/8-1:0] m_axis_bramio_61_tkeep,
    output [C_INOUT_BRAM_61_DMWIDTH/8-1:0] m_axis_bramio_61_tstrb,
    output [C_INOUT_BRAM_61_DMWIDTH-1:0] m_axis_bramio_61_tdata,
    input m_axis_bramio_61_tready,
    //in-out BRAM AXI-Stream output interface 62
    output m_axis_bramio_62_tlast,
    output m_axis_bramio_62_tvalid,
    output [C_INOUT_BRAM_62_DMWIDTH/8-1:0] m_axis_bramio_62_tkeep,
    output [C_INOUT_BRAM_62_DMWIDTH/8-1:0] m_axis_bramio_62_tstrb,
    output [C_INOUT_BRAM_62_DMWIDTH-1:0] m_axis_bramio_62_tdata,
    input m_axis_bramio_62_tready,
    //in-out BRAM AXI-Stream output interface 63
    output m_axis_bramio_63_tlast,
    output m_axis_bramio_63_tvalid,
    output [C_INOUT_BRAM_63_DMWIDTH/8-1:0] m_axis_bramio_63_tkeep,
    output [C_INOUT_BRAM_63_DMWIDTH/8-1:0] m_axis_bramio_63_tstrb,
    output [C_INOUT_BRAM_63_DMWIDTH-1:0] m_axis_bramio_63_tdata,
    input m_axis_bramio_63_tready,
    //in-out BRAM AXI-Stream output interface 64
    output m_axis_bramio_64_tlast,
    output m_axis_bramio_64_tvalid,
    output [C_INOUT_BRAM_64_DMWIDTH/8-1:0] m_axis_bramio_64_tkeep,
    output [C_INOUT_BRAM_64_DMWIDTH/8-1:0] m_axis_bramio_64_tstrb,
    output [C_INOUT_BRAM_64_DMWIDTH-1:0] m_axis_bramio_64_tdata,
    input m_axis_bramio_64_tready,
    //in-out BRAM AXI-Stream output interface 65
    output m_axis_bramio_65_tlast,
    output m_axis_bramio_65_tvalid,
    output [C_INOUT_BRAM_65_DMWIDTH/8-1:0] m_axis_bramio_65_tkeep,
    output [C_INOUT_BRAM_65_DMWIDTH/8-1:0] m_axis_bramio_65_tstrb,
    output [C_INOUT_BRAM_65_DMWIDTH-1:0] m_axis_bramio_65_tdata,
    input m_axis_bramio_65_tready,
    //in-out BRAM AXI-Stream output interface 66
    output m_axis_bramio_66_tlast,
    output m_axis_bramio_66_tvalid,
    output [C_INOUT_BRAM_66_DMWIDTH/8-1:0] m_axis_bramio_66_tkeep,
    output [C_INOUT_BRAM_66_DMWIDTH/8-1:0] m_axis_bramio_66_tstrb,
    output [C_INOUT_BRAM_66_DMWIDTH-1:0] m_axis_bramio_66_tdata,
    input m_axis_bramio_66_tready,
    //in-out BRAM AXI-Stream output interface 67
    output m_axis_bramio_67_tlast,
    output m_axis_bramio_67_tvalid,
    output [C_INOUT_BRAM_67_DMWIDTH/8-1:0] m_axis_bramio_67_tkeep,
    output [C_INOUT_BRAM_67_DMWIDTH/8-1:0] m_axis_bramio_67_tstrb,
    output [C_INOUT_BRAM_67_DMWIDTH-1:0] m_axis_bramio_67_tdata,
    input m_axis_bramio_67_tready,
    //in-out BRAM AXI-Stream output interface 68
    output m_axis_bramio_68_tlast,
    output m_axis_bramio_68_tvalid,
    output [C_INOUT_BRAM_68_DMWIDTH/8-1:0] m_axis_bramio_68_tkeep,
    output [C_INOUT_BRAM_68_DMWIDTH/8-1:0] m_axis_bramio_68_tstrb,
    output [C_INOUT_BRAM_68_DMWIDTH-1:0] m_axis_bramio_68_tdata,
    input m_axis_bramio_68_tready,
    //in-out BRAM AXI-Stream output interface 69
    output m_axis_bramio_69_tlast,
    output m_axis_bramio_69_tvalid,
    output [C_INOUT_BRAM_69_DMWIDTH/8-1:0] m_axis_bramio_69_tkeep,
    output [C_INOUT_BRAM_69_DMWIDTH/8-1:0] m_axis_bramio_69_tstrb,
    output [C_INOUT_BRAM_69_DMWIDTH-1:0] m_axis_bramio_69_tdata,
    input m_axis_bramio_69_tready,
    //in-out BRAM AXI-Stream output interface 70
    output m_axis_bramio_70_tlast,
    output m_axis_bramio_70_tvalid,
    output [C_INOUT_BRAM_70_DMWIDTH/8-1:0] m_axis_bramio_70_tkeep,
    output [C_INOUT_BRAM_70_DMWIDTH/8-1:0] m_axis_bramio_70_tstrb,
    output [C_INOUT_BRAM_70_DMWIDTH-1:0] m_axis_bramio_70_tdata,
    input m_axis_bramio_70_tready,
    //in-out BRAM AXI-Stream output interface 71
    output m_axis_bramio_71_tlast,
    output m_axis_bramio_71_tvalid,
    output [C_INOUT_BRAM_71_DMWIDTH/8-1:0] m_axis_bramio_71_tkeep,
    output [C_INOUT_BRAM_71_DMWIDTH/8-1:0] m_axis_bramio_71_tstrb,
    output [C_INOUT_BRAM_71_DMWIDTH-1:0] m_axis_bramio_71_tdata,
    input m_axis_bramio_71_tready,
    //in-out BRAM AXI-Stream output interface 72
    output m_axis_bramio_72_tlast,
    output m_axis_bramio_72_tvalid,
    output [C_INOUT_BRAM_72_DMWIDTH/8-1:0] m_axis_bramio_72_tkeep,
    output [C_INOUT_BRAM_72_DMWIDTH/8-1:0] m_axis_bramio_72_tstrb,
    output [C_INOUT_BRAM_72_DMWIDTH-1:0] m_axis_bramio_72_tdata,
    input m_axis_bramio_72_tready,
    //in-out BRAM AXI-Stream output interface 73
    output m_axis_bramio_73_tlast,
    output m_axis_bramio_73_tvalid,
    output [C_INOUT_BRAM_73_DMWIDTH/8-1:0] m_axis_bramio_73_tkeep,
    output [C_INOUT_BRAM_73_DMWIDTH/8-1:0] m_axis_bramio_73_tstrb,
    output [C_INOUT_BRAM_73_DMWIDTH-1:0] m_axis_bramio_73_tdata,
    input m_axis_bramio_73_tready,
    //in-out BRAM AXI-Stream output interface 74
    output m_axis_bramio_74_tlast,
    output m_axis_bramio_74_tvalid,
    output [C_INOUT_BRAM_74_DMWIDTH/8-1:0] m_axis_bramio_74_tkeep,
    output [C_INOUT_BRAM_74_DMWIDTH/8-1:0] m_axis_bramio_74_tstrb,
    output [C_INOUT_BRAM_74_DMWIDTH-1:0] m_axis_bramio_74_tdata,
    input m_axis_bramio_74_tready,
    //in-out BRAM AXI-Stream output interface 75
    output m_axis_bramio_75_tlast,
    output m_axis_bramio_75_tvalid,
    output [C_INOUT_BRAM_75_DMWIDTH/8-1:0] m_axis_bramio_75_tkeep,
    output [C_INOUT_BRAM_75_DMWIDTH/8-1:0] m_axis_bramio_75_tstrb,
    output [C_INOUT_BRAM_75_DMWIDTH-1:0] m_axis_bramio_75_tdata,
    input m_axis_bramio_75_tready,
    //in-out BRAM AXI-Stream output interface 76
    output m_axis_bramio_76_tlast,
    output m_axis_bramio_76_tvalid,
    output [C_INOUT_BRAM_76_DMWIDTH/8-1:0] m_axis_bramio_76_tkeep,
    output [C_INOUT_BRAM_76_DMWIDTH/8-1:0] m_axis_bramio_76_tstrb,
    output [C_INOUT_BRAM_76_DMWIDTH-1:0] m_axis_bramio_76_tdata,
    input m_axis_bramio_76_tready,
    //in-out BRAM AXI-Stream output interface 77
    output m_axis_bramio_77_tlast,
    output m_axis_bramio_77_tvalid,
    output [C_INOUT_BRAM_77_DMWIDTH/8-1:0] m_axis_bramio_77_tkeep,
    output [C_INOUT_BRAM_77_DMWIDTH/8-1:0] m_axis_bramio_77_tstrb,
    output [C_INOUT_BRAM_77_DMWIDTH-1:0] m_axis_bramio_77_tdata,
    input m_axis_bramio_77_tready,
    //in-out BRAM AXI-Stream output interface 78
    output m_axis_bramio_78_tlast,
    output m_axis_bramio_78_tvalid,
    output [C_INOUT_BRAM_78_DMWIDTH/8-1:0] m_axis_bramio_78_tkeep,
    output [C_INOUT_BRAM_78_DMWIDTH/8-1:0] m_axis_bramio_78_tstrb,
    output [C_INOUT_BRAM_78_DMWIDTH-1:0] m_axis_bramio_78_tdata,
    input m_axis_bramio_78_tready,
    //in-out BRAM AXI-Stream output interface 79
    output m_axis_bramio_79_tlast,
    output m_axis_bramio_79_tvalid,
    output [C_INOUT_BRAM_79_DMWIDTH/8-1:0] m_axis_bramio_79_tkeep,
    output [C_INOUT_BRAM_79_DMWIDTH/8-1:0] m_axis_bramio_79_tstrb,
    output [C_INOUT_BRAM_79_DMWIDTH-1:0] m_axis_bramio_79_tdata,
    input m_axis_bramio_79_tready,
    //in-out BRAM AXI-Stream output interface 80
    output m_axis_bramio_80_tlast,
    output m_axis_bramio_80_tvalid,
    output [C_INOUT_BRAM_80_DMWIDTH/8-1:0] m_axis_bramio_80_tkeep,
    output [C_INOUT_BRAM_80_DMWIDTH/8-1:0] m_axis_bramio_80_tstrb,
    output [C_INOUT_BRAM_80_DMWIDTH-1:0] m_axis_bramio_80_tdata,
    input m_axis_bramio_80_tready,
    //in-out BRAM AXI-Stream output interface 81
    output m_axis_bramio_81_tlast,
    output m_axis_bramio_81_tvalid,
    output [C_INOUT_BRAM_81_DMWIDTH/8-1:0] m_axis_bramio_81_tkeep,
    output [C_INOUT_BRAM_81_DMWIDTH/8-1:0] m_axis_bramio_81_tstrb,
    output [C_INOUT_BRAM_81_DMWIDTH-1:0] m_axis_bramio_81_tdata,
    input m_axis_bramio_81_tready,
    //in-out BRAM AXI-Stream output interface 82
    output m_axis_bramio_82_tlast,
    output m_axis_bramio_82_tvalid,
    output [C_INOUT_BRAM_82_DMWIDTH/8-1:0] m_axis_bramio_82_tkeep,
    output [C_INOUT_BRAM_82_DMWIDTH/8-1:0] m_axis_bramio_82_tstrb,
    output [C_INOUT_BRAM_82_DMWIDTH-1:0] m_axis_bramio_82_tdata,
    input m_axis_bramio_82_tready,
    //in-out BRAM AXI-Stream output interface 83
    output m_axis_bramio_83_tlast,
    output m_axis_bramio_83_tvalid,
    output [C_INOUT_BRAM_83_DMWIDTH/8-1:0] m_axis_bramio_83_tkeep,
    output [C_INOUT_BRAM_83_DMWIDTH/8-1:0] m_axis_bramio_83_tstrb,
    output [C_INOUT_BRAM_83_DMWIDTH-1:0] m_axis_bramio_83_tdata,
    input m_axis_bramio_83_tready,
    //in-out BRAM AXI-Stream output interface 84
    output m_axis_bramio_84_tlast,
    output m_axis_bramio_84_tvalid,
    output [C_INOUT_BRAM_84_DMWIDTH/8-1:0] m_axis_bramio_84_tkeep,
    output [C_INOUT_BRAM_84_DMWIDTH/8-1:0] m_axis_bramio_84_tstrb,
    output [C_INOUT_BRAM_84_DMWIDTH-1:0] m_axis_bramio_84_tdata,
    input m_axis_bramio_84_tready,
    //in-out BRAM AXI-Stream output interface 85
    output m_axis_bramio_85_tlast,
    output m_axis_bramio_85_tvalid,
    output [C_INOUT_BRAM_85_DMWIDTH/8-1:0] m_axis_bramio_85_tkeep,
    output [C_INOUT_BRAM_85_DMWIDTH/8-1:0] m_axis_bramio_85_tstrb,
    output [C_INOUT_BRAM_85_DMWIDTH-1:0] m_axis_bramio_85_tdata,
    input m_axis_bramio_85_tready,
    //in-out BRAM AXI-Stream output interface 86
    output m_axis_bramio_86_tlast,
    output m_axis_bramio_86_tvalid,
    output [C_INOUT_BRAM_86_DMWIDTH/8-1:0] m_axis_bramio_86_tkeep,
    output [C_INOUT_BRAM_86_DMWIDTH/8-1:0] m_axis_bramio_86_tstrb,
    output [C_INOUT_BRAM_86_DMWIDTH-1:0] m_axis_bramio_86_tdata,
    input m_axis_bramio_86_tready,
    //in-out BRAM AXI-Stream output interface 87
    output m_axis_bramio_87_tlast,
    output m_axis_bramio_87_tvalid,
    output [C_INOUT_BRAM_87_DMWIDTH/8-1:0] m_axis_bramio_87_tkeep,
    output [C_INOUT_BRAM_87_DMWIDTH/8-1:0] m_axis_bramio_87_tstrb,
    output [C_INOUT_BRAM_87_DMWIDTH-1:0] m_axis_bramio_87_tdata,
    input m_axis_bramio_87_tready,
    //in-out BRAM AXI-Stream output interface 88
    output m_axis_bramio_88_tlast,
    output m_axis_bramio_88_tvalid,
    output [C_INOUT_BRAM_88_DMWIDTH/8-1:0] m_axis_bramio_88_tkeep,
    output [C_INOUT_BRAM_88_DMWIDTH/8-1:0] m_axis_bramio_88_tstrb,
    output [C_INOUT_BRAM_88_DMWIDTH-1:0] m_axis_bramio_88_tdata,
    input m_axis_bramio_88_tready,
    //in-out BRAM AXI-Stream output interface 89
    output m_axis_bramio_89_tlast,
    output m_axis_bramio_89_tvalid,
    output [C_INOUT_BRAM_89_DMWIDTH/8-1:0] m_axis_bramio_89_tkeep,
    output [C_INOUT_BRAM_89_DMWIDTH/8-1:0] m_axis_bramio_89_tstrb,
    output [C_INOUT_BRAM_89_DMWIDTH-1:0] m_axis_bramio_89_tdata,
    input m_axis_bramio_89_tready,
    //in-out BRAM AXI-Stream output interface 90
    output m_axis_bramio_90_tlast,
    output m_axis_bramio_90_tvalid,
    output [C_INOUT_BRAM_90_DMWIDTH/8-1:0] m_axis_bramio_90_tkeep,
    output [C_INOUT_BRAM_90_DMWIDTH/8-1:0] m_axis_bramio_90_tstrb,
    output [C_INOUT_BRAM_90_DMWIDTH-1:0] m_axis_bramio_90_tdata,
    input m_axis_bramio_90_tready,
    //in-out BRAM AXI-Stream output interface 91
    output m_axis_bramio_91_tlast,
    output m_axis_bramio_91_tvalid,
    output [C_INOUT_BRAM_91_DMWIDTH/8-1:0] m_axis_bramio_91_tkeep,
    output [C_INOUT_BRAM_91_DMWIDTH/8-1:0] m_axis_bramio_91_tstrb,
    output [C_INOUT_BRAM_91_DMWIDTH-1:0] m_axis_bramio_91_tdata,
    input m_axis_bramio_91_tready,
    //in-out BRAM AXI-Stream output interface 92
    output m_axis_bramio_92_tlast,
    output m_axis_bramio_92_tvalid,
    output [C_INOUT_BRAM_92_DMWIDTH/8-1:0] m_axis_bramio_92_tkeep,
    output [C_INOUT_BRAM_92_DMWIDTH/8-1:0] m_axis_bramio_92_tstrb,
    output [C_INOUT_BRAM_92_DMWIDTH-1:0] m_axis_bramio_92_tdata,
    input m_axis_bramio_92_tready,
    //in-out BRAM AXI-Stream output interface 93
    output m_axis_bramio_93_tlast,
    output m_axis_bramio_93_tvalid,
    output [C_INOUT_BRAM_93_DMWIDTH/8-1:0] m_axis_bramio_93_tkeep,
    output [C_INOUT_BRAM_93_DMWIDTH/8-1:0] m_axis_bramio_93_tstrb,
    output [C_INOUT_BRAM_93_DMWIDTH-1:0] m_axis_bramio_93_tdata,
    input m_axis_bramio_93_tready,
    //in-out BRAM AXI-Stream output interface 94
    output m_axis_bramio_94_tlast,
    output m_axis_bramio_94_tvalid,
    output [C_INOUT_BRAM_94_DMWIDTH/8-1:0] m_axis_bramio_94_tkeep,
    output [C_INOUT_BRAM_94_DMWIDTH/8-1:0] m_axis_bramio_94_tstrb,
    output [C_INOUT_BRAM_94_DMWIDTH-1:0] m_axis_bramio_94_tdata,
    input m_axis_bramio_94_tready,
    //in-out BRAM AXI-Stream output interface 95
    output m_axis_bramio_95_tlast,
    output m_axis_bramio_95_tvalid,
    output [C_INOUT_BRAM_95_DMWIDTH/8-1:0] m_axis_bramio_95_tkeep,
    output [C_INOUT_BRAM_95_DMWIDTH/8-1:0] m_axis_bramio_95_tstrb,
    output [C_INOUT_BRAM_95_DMWIDTH-1:0] m_axis_bramio_95_tdata,
    input m_axis_bramio_95_tready,
    //in-out BRAM AXI-Stream output interface 96
    output m_axis_bramio_96_tlast,
    output m_axis_bramio_96_tvalid,
    output [C_INOUT_BRAM_96_DMWIDTH/8-1:0] m_axis_bramio_96_tkeep,
    output [C_INOUT_BRAM_96_DMWIDTH/8-1:0] m_axis_bramio_96_tstrb,
    output [C_INOUT_BRAM_96_DMWIDTH-1:0] m_axis_bramio_96_tdata,
    input m_axis_bramio_96_tready,
    //in-out BRAM AXI-Stream output interface 97
    output m_axis_bramio_97_tlast,
    output m_axis_bramio_97_tvalid,
    output [C_INOUT_BRAM_97_DMWIDTH/8-1:0] m_axis_bramio_97_tkeep,
    output [C_INOUT_BRAM_97_DMWIDTH/8-1:0] m_axis_bramio_97_tstrb,
    output [C_INOUT_BRAM_97_DMWIDTH-1:0] m_axis_bramio_97_tdata,
    input m_axis_bramio_97_tready,
    //in-out BRAM AXI-Stream output interface 98
    output m_axis_bramio_98_tlast,
    output m_axis_bramio_98_tvalid,
    output [C_INOUT_BRAM_98_DMWIDTH/8-1:0] m_axis_bramio_98_tkeep,
    output [C_INOUT_BRAM_98_DMWIDTH/8-1:0] m_axis_bramio_98_tstrb,
    output [C_INOUT_BRAM_98_DMWIDTH-1:0] m_axis_bramio_98_tdata,
    input m_axis_bramio_98_tready,
    //in-out BRAM AXI-Stream output interface 99
    output m_axis_bramio_99_tlast,
    output m_axis_bramio_99_tvalid,
    output [C_INOUT_BRAM_99_DMWIDTH/8-1:0] m_axis_bramio_99_tkeep,
    output [C_INOUT_BRAM_99_DMWIDTH/8-1:0] m_axis_bramio_99_tstrb,
    output [C_INOUT_BRAM_99_DMWIDTH-1:0] m_axis_bramio_99_tdata,
    input m_axis_bramio_99_tready,
    //in-out BRAM AXI-Stream output interface 100
    output m_axis_bramio_100_tlast,
    output m_axis_bramio_100_tvalid,
    output [C_INOUT_BRAM_100_DMWIDTH/8-1:0] m_axis_bramio_100_tkeep,
    output [C_INOUT_BRAM_100_DMWIDTH/8-1:0] m_axis_bramio_100_tstrb,
    output [C_INOUT_BRAM_100_DMWIDTH-1:0] m_axis_bramio_100_tdata,
    input m_axis_bramio_100_tready,
    //in-out BRAM AXI-Stream output interface 101
    output m_axis_bramio_101_tlast,
    output m_axis_bramio_101_tvalid,
    output [C_INOUT_BRAM_101_DMWIDTH/8-1:0] m_axis_bramio_101_tkeep,
    output [C_INOUT_BRAM_101_DMWIDTH/8-1:0] m_axis_bramio_101_tstrb,
    output [C_INOUT_BRAM_101_DMWIDTH-1:0] m_axis_bramio_101_tdata,
    input m_axis_bramio_101_tready,
    //in-out BRAM AXI-Stream output interface 102
    output m_axis_bramio_102_tlast,
    output m_axis_bramio_102_tvalid,
    output [C_INOUT_BRAM_102_DMWIDTH/8-1:0] m_axis_bramio_102_tkeep,
    output [C_INOUT_BRAM_102_DMWIDTH/8-1:0] m_axis_bramio_102_tstrb,
    output [C_INOUT_BRAM_102_DMWIDTH-1:0] m_axis_bramio_102_tdata,
    input m_axis_bramio_102_tready,
    //in-out BRAM AXI-Stream output interface 103
    output m_axis_bramio_103_tlast,
    output m_axis_bramio_103_tvalid,
    output [C_INOUT_BRAM_103_DMWIDTH/8-1:0] m_axis_bramio_103_tkeep,
    output [C_INOUT_BRAM_103_DMWIDTH/8-1:0] m_axis_bramio_103_tstrb,
    output [C_INOUT_BRAM_103_DMWIDTH-1:0] m_axis_bramio_103_tdata,
    input m_axis_bramio_103_tready,
    //in-out BRAM AXI-Stream output interface 104
    output m_axis_bramio_104_tlast,
    output m_axis_bramio_104_tvalid,
    output [C_INOUT_BRAM_104_DMWIDTH/8-1:0] m_axis_bramio_104_tkeep,
    output [C_INOUT_BRAM_104_DMWIDTH/8-1:0] m_axis_bramio_104_tstrb,
    output [C_INOUT_BRAM_104_DMWIDTH-1:0] m_axis_bramio_104_tdata,
    input m_axis_bramio_104_tready,
    //in-out BRAM AXI-Stream output interface 105
    output m_axis_bramio_105_tlast,
    output m_axis_bramio_105_tvalid,
    output [C_INOUT_BRAM_105_DMWIDTH/8-1:0] m_axis_bramio_105_tkeep,
    output [C_INOUT_BRAM_105_DMWIDTH/8-1:0] m_axis_bramio_105_tstrb,
    output [C_INOUT_BRAM_105_DMWIDTH-1:0] m_axis_bramio_105_tdata,
    input m_axis_bramio_105_tready,
    //in-out BRAM AXI-Stream output interface 106
    output m_axis_bramio_106_tlast,
    output m_axis_bramio_106_tvalid,
    output [C_INOUT_BRAM_106_DMWIDTH/8-1:0] m_axis_bramio_106_tkeep,
    output [C_INOUT_BRAM_106_DMWIDTH/8-1:0] m_axis_bramio_106_tstrb,
    output [C_INOUT_BRAM_106_DMWIDTH-1:0] m_axis_bramio_106_tdata,
    input m_axis_bramio_106_tready,
    //in-out BRAM AXI-Stream output interface 107
    output m_axis_bramio_107_tlast,
    output m_axis_bramio_107_tvalid,
    output [C_INOUT_BRAM_107_DMWIDTH/8-1:0] m_axis_bramio_107_tkeep,
    output [C_INOUT_BRAM_107_DMWIDTH/8-1:0] m_axis_bramio_107_tstrb,
    output [C_INOUT_BRAM_107_DMWIDTH-1:0] m_axis_bramio_107_tdata,
    input m_axis_bramio_107_tready,
    //in-out BRAM AXI-Stream output interface 108
    output m_axis_bramio_108_tlast,
    output m_axis_bramio_108_tvalid,
    output [C_INOUT_BRAM_108_DMWIDTH/8-1:0] m_axis_bramio_108_tkeep,
    output [C_INOUT_BRAM_108_DMWIDTH/8-1:0] m_axis_bramio_108_tstrb,
    output [C_INOUT_BRAM_108_DMWIDTH-1:0] m_axis_bramio_108_tdata,
    input m_axis_bramio_108_tready,
    //in-out BRAM AXI-Stream output interface 109
    output m_axis_bramio_109_tlast,
    output m_axis_bramio_109_tvalid,
    output [C_INOUT_BRAM_109_DMWIDTH/8-1:0] m_axis_bramio_109_tkeep,
    output [C_INOUT_BRAM_109_DMWIDTH/8-1:0] m_axis_bramio_109_tstrb,
    output [C_INOUT_BRAM_109_DMWIDTH-1:0] m_axis_bramio_109_tdata,
    input m_axis_bramio_109_tready,
    //in-out BRAM AXI-Stream output interface 110
    output m_axis_bramio_110_tlast,
    output m_axis_bramio_110_tvalid,
    output [C_INOUT_BRAM_110_DMWIDTH/8-1:0] m_axis_bramio_110_tkeep,
    output [C_INOUT_BRAM_110_DMWIDTH/8-1:0] m_axis_bramio_110_tstrb,
    output [C_INOUT_BRAM_110_DMWIDTH-1:0] m_axis_bramio_110_tdata,
    input m_axis_bramio_110_tready,
    //in-out BRAM AXI-Stream output interface 111
    output m_axis_bramio_111_tlast,
    output m_axis_bramio_111_tvalid,
    output [C_INOUT_BRAM_111_DMWIDTH/8-1:0] m_axis_bramio_111_tkeep,
    output [C_INOUT_BRAM_111_DMWIDTH/8-1:0] m_axis_bramio_111_tstrb,
    output [C_INOUT_BRAM_111_DMWIDTH-1:0] m_axis_bramio_111_tdata,
    input m_axis_bramio_111_tready,
    //in-out BRAM AXI-Stream output interface 112
    output m_axis_bramio_112_tlast,
    output m_axis_bramio_112_tvalid,
    output [C_INOUT_BRAM_112_DMWIDTH/8-1:0] m_axis_bramio_112_tkeep,
    output [C_INOUT_BRAM_112_DMWIDTH/8-1:0] m_axis_bramio_112_tstrb,
    output [C_INOUT_BRAM_112_DMWIDTH-1:0] m_axis_bramio_112_tdata,
    input m_axis_bramio_112_tready,
    //in-out BRAM AXI-Stream output interface 113
    output m_axis_bramio_113_tlast,
    output m_axis_bramio_113_tvalid,
    output [C_INOUT_BRAM_113_DMWIDTH/8-1:0] m_axis_bramio_113_tkeep,
    output [C_INOUT_BRAM_113_DMWIDTH/8-1:0] m_axis_bramio_113_tstrb,
    output [C_INOUT_BRAM_113_DMWIDTH-1:0] m_axis_bramio_113_tdata,
    input m_axis_bramio_113_tready,
    //in-out BRAM AXI-Stream output interface 114
    output m_axis_bramio_114_tlast,
    output m_axis_bramio_114_tvalid,
    output [C_INOUT_BRAM_114_DMWIDTH/8-1:0] m_axis_bramio_114_tkeep,
    output [C_INOUT_BRAM_114_DMWIDTH/8-1:0] m_axis_bramio_114_tstrb,
    output [C_INOUT_BRAM_114_DMWIDTH-1:0] m_axis_bramio_114_tdata,
    input m_axis_bramio_114_tready,
    //in-out BRAM AXI-Stream output interface 115
    output m_axis_bramio_115_tlast,
    output m_axis_bramio_115_tvalid,
    output [C_INOUT_BRAM_115_DMWIDTH/8-1:0] m_axis_bramio_115_tkeep,
    output [C_INOUT_BRAM_115_DMWIDTH/8-1:0] m_axis_bramio_115_tstrb,
    output [C_INOUT_BRAM_115_DMWIDTH-1:0] m_axis_bramio_115_tdata,
    input m_axis_bramio_115_tready,
    //in-out BRAM AXI-Stream output interface 116
    output m_axis_bramio_116_tlast,
    output m_axis_bramio_116_tvalid,
    output [C_INOUT_BRAM_116_DMWIDTH/8-1:0] m_axis_bramio_116_tkeep,
    output [C_INOUT_BRAM_116_DMWIDTH/8-1:0] m_axis_bramio_116_tstrb,
    output [C_INOUT_BRAM_116_DMWIDTH-1:0] m_axis_bramio_116_tdata,
    input m_axis_bramio_116_tready,
    //in-out BRAM AXI-Stream output interface 117
    output m_axis_bramio_117_tlast,
    output m_axis_bramio_117_tvalid,
    output [C_INOUT_BRAM_117_DMWIDTH/8-1:0] m_axis_bramio_117_tkeep,
    output [C_INOUT_BRAM_117_DMWIDTH/8-1:0] m_axis_bramio_117_tstrb,
    output [C_INOUT_BRAM_117_DMWIDTH-1:0] m_axis_bramio_117_tdata,
    input m_axis_bramio_117_tready,
    //in-out BRAM AXI-Stream output interface 118
    output m_axis_bramio_118_tlast,
    output m_axis_bramio_118_tvalid,
    output [C_INOUT_BRAM_118_DMWIDTH/8-1:0] m_axis_bramio_118_tkeep,
    output [C_INOUT_BRAM_118_DMWIDTH/8-1:0] m_axis_bramio_118_tstrb,
    output [C_INOUT_BRAM_118_DMWIDTH-1:0] m_axis_bramio_118_tdata,
    input m_axis_bramio_118_tready,
    //in-out BRAM AXI-Stream output interface 119
    output m_axis_bramio_119_tlast,
    output m_axis_bramio_119_tvalid,
    output [C_INOUT_BRAM_119_DMWIDTH/8-1:0] m_axis_bramio_119_tkeep,
    output [C_INOUT_BRAM_119_DMWIDTH/8-1:0] m_axis_bramio_119_tstrb,
    output [C_INOUT_BRAM_119_DMWIDTH-1:0] m_axis_bramio_119_tdata,
    input m_axis_bramio_119_tready,
    //in-out BRAM AXI-Stream output interface 120
    output m_axis_bramio_120_tlast,
    output m_axis_bramio_120_tvalid,
    output [C_INOUT_BRAM_120_DMWIDTH/8-1:0] m_axis_bramio_120_tkeep,
    output [C_INOUT_BRAM_120_DMWIDTH/8-1:0] m_axis_bramio_120_tstrb,
    output [C_INOUT_BRAM_120_DMWIDTH-1:0] m_axis_bramio_120_tdata,
    input m_axis_bramio_120_tready,
    //in-out BRAM AXI-Stream output interface 121
    output m_axis_bramio_121_tlast,
    output m_axis_bramio_121_tvalid,
    output [C_INOUT_BRAM_121_DMWIDTH/8-1:0] m_axis_bramio_121_tkeep,
    output [C_INOUT_BRAM_121_DMWIDTH/8-1:0] m_axis_bramio_121_tstrb,
    output [C_INOUT_BRAM_121_DMWIDTH-1:0] m_axis_bramio_121_tdata,
    input m_axis_bramio_121_tready,
    //in-out BRAM AXI-Stream output interface 122
    output m_axis_bramio_122_tlast,
    output m_axis_bramio_122_tvalid,
    output [C_INOUT_BRAM_122_DMWIDTH/8-1:0] m_axis_bramio_122_tkeep,
    output [C_INOUT_BRAM_122_DMWIDTH/8-1:0] m_axis_bramio_122_tstrb,
    output [C_INOUT_BRAM_122_DMWIDTH-1:0] m_axis_bramio_122_tdata,
    input m_axis_bramio_122_tready,
    //in-out BRAM AXI-Stream output interface 123
    output m_axis_bramio_123_tlast,
    output m_axis_bramio_123_tvalid,
    output [C_INOUT_BRAM_123_DMWIDTH/8-1:0] m_axis_bramio_123_tkeep,
    output [C_INOUT_BRAM_123_DMWIDTH/8-1:0] m_axis_bramio_123_tstrb,
    output [C_INOUT_BRAM_123_DMWIDTH-1:0] m_axis_bramio_123_tdata,
    input m_axis_bramio_123_tready,
    //in-out BRAM AXI-Stream output interface 124
    output m_axis_bramio_124_tlast,
    output m_axis_bramio_124_tvalid,
    output [C_INOUT_BRAM_124_DMWIDTH/8-1:0] m_axis_bramio_124_tkeep,
    output [C_INOUT_BRAM_124_DMWIDTH/8-1:0] m_axis_bramio_124_tstrb,
    output [C_INOUT_BRAM_124_DMWIDTH-1:0] m_axis_bramio_124_tdata,
    input m_axis_bramio_124_tready,
    //in-out BRAM AXI-Stream output interface 125
    output m_axis_bramio_125_tlast,
    output m_axis_bramio_125_tvalid,
    output [C_INOUT_BRAM_125_DMWIDTH/8-1:0] m_axis_bramio_125_tkeep,
    output [C_INOUT_BRAM_125_DMWIDTH/8-1:0] m_axis_bramio_125_tstrb,
    output [C_INOUT_BRAM_125_DMWIDTH-1:0] m_axis_bramio_125_tdata,
    input m_axis_bramio_125_tready,
    //in-out BRAM AXI-Stream output interface 126
    output m_axis_bramio_126_tlast,
    output m_axis_bramio_126_tvalid,
    output [C_INOUT_BRAM_126_DMWIDTH/8-1:0] m_axis_bramio_126_tkeep,
    output [C_INOUT_BRAM_126_DMWIDTH/8-1:0] m_axis_bramio_126_tstrb,
    output [C_INOUT_BRAM_126_DMWIDTH-1:0] m_axis_bramio_126_tdata,
    input m_axis_bramio_126_tready,
    //in-out BRAM AXI-Stream output interface 127
    output m_axis_bramio_127_tlast,
    output m_axis_bramio_127_tvalid,
    output [C_INOUT_BRAM_127_DMWIDTH/8-1:0] m_axis_bramio_127_tkeep,
    output [C_INOUT_BRAM_127_DMWIDTH/8-1:0] m_axis_bramio_127_tstrb,
    output [C_INOUT_BRAM_127_DMWIDTH-1:0] m_axis_bramio_127_tdata,
    input m_axis_bramio_127_tready,
    //-----------------------------------------------------------
    //out AXI-Stream output interface 0
    output m_axis_bram_0_tlast,
    output m_axis_bram_0_tvalid,
    output [C_OUTPUT_BRAM_0_DMWIDTH/8-1:0] m_axis_bram_0_tkeep,
    output [C_OUTPUT_BRAM_0_DMWIDTH/8-1:0] m_axis_bram_0_tstrb,
    output [C_OUTPUT_BRAM_0_DMWIDTH-1:0] m_axis_bram_0_tdata,
    input m_axis_bram_0_tready,
    input [C_OUTPUT_BRAM_0_ADDR_WIDTH-1:0] ap_bram_oarg_0_addr0,
    input [C_OUTPUT_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_din0,
    output [C_OUTPUT_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_dout0,
    input ap_bram_oarg_0_clk0,
    input ap_bram_oarg_0_rst0,
    input [C_OUTPUT_BRAM_0_WIDTH/8-1:0] ap_bram_oarg_0_we0,
    input ap_bram_oarg_0_en0,
    input [C_OUTPUT_BRAM_0_ADDR_WIDTH-1:0] ap_bram_oarg_0_addr1,
    input [C_OUTPUT_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_din1,
    output [C_OUTPUT_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_dout1,
    input ap_bram_oarg_0_clk1,
    input ap_bram_oarg_0_rst1,
    input [C_OUTPUT_BRAM_0_WIDTH/8-1:0] ap_bram_oarg_0_we1,
    input ap_bram_oarg_0_en1,
    //out AXI-Stream output interface 1
    output m_axis_bram_1_tlast,
    output m_axis_bram_1_tvalid,
    output [C_OUTPUT_BRAM_1_DMWIDTH/8-1:0] m_axis_bram_1_tkeep,
    output [C_OUTPUT_BRAM_1_DMWIDTH/8-1:0] m_axis_bram_1_tstrb,
    output [C_OUTPUT_BRAM_1_DMWIDTH-1:0] m_axis_bram_1_tdata,
    input m_axis_bram_1_tready,
    input [C_OUTPUT_BRAM_1_ADDR_WIDTH-1:0] ap_bram_oarg_1_addr0,
    input [C_OUTPUT_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_din0,
    output [C_OUTPUT_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_dout0,
    input ap_bram_oarg_1_clk0,
    input ap_bram_oarg_1_rst0,
    input [C_OUTPUT_BRAM_1_WIDTH/8-1:0] ap_bram_oarg_1_we0,
    input ap_bram_oarg_1_en0,
    input [C_OUTPUT_BRAM_1_ADDR_WIDTH-1:0] ap_bram_oarg_1_addr1,
    input [C_OUTPUT_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_din1,
    output [C_OUTPUT_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_dout1,
    input ap_bram_oarg_1_clk1,
    input ap_bram_oarg_1_rst1,
    input [C_OUTPUT_BRAM_1_WIDTH/8-1:0] ap_bram_oarg_1_we1,
    input ap_bram_oarg_1_en1,
    //out AXI-Stream output interface 2
    output m_axis_bram_2_tlast,
    output m_axis_bram_2_tvalid,
    output [C_OUTPUT_BRAM_2_DMWIDTH/8-1:0] m_axis_bram_2_tkeep,
    output [C_OUTPUT_BRAM_2_DMWIDTH/8-1:0] m_axis_bram_2_tstrb,
    output [C_OUTPUT_BRAM_2_DMWIDTH-1:0] m_axis_bram_2_tdata,
    input m_axis_bram_2_tready,
    input [C_OUTPUT_BRAM_2_ADDR_WIDTH-1:0] ap_bram_oarg_2_addr0,
    input [C_OUTPUT_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_din0,
    output [C_OUTPUT_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_dout0,
    input ap_bram_oarg_2_clk0,
    input ap_bram_oarg_2_rst0,
    input [C_OUTPUT_BRAM_2_WIDTH/8-1:0] ap_bram_oarg_2_we0,
    input ap_bram_oarg_2_en0,
    input [C_OUTPUT_BRAM_2_ADDR_WIDTH-1:0] ap_bram_oarg_2_addr1,
    input [C_OUTPUT_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_din1,
    output [C_OUTPUT_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_dout1,
    input ap_bram_oarg_2_clk1,
    input ap_bram_oarg_2_rst1,
    input [C_OUTPUT_BRAM_2_WIDTH/8-1:0] ap_bram_oarg_2_we1,
    input ap_bram_oarg_2_en1,
    //out AXI-Stream output interface 3
    output m_axis_bram_3_tlast,
    output m_axis_bram_3_tvalid,
    output [C_OUTPUT_BRAM_3_DMWIDTH/8-1:0] m_axis_bram_3_tkeep,
    output [C_OUTPUT_BRAM_3_DMWIDTH/8-1:0] m_axis_bram_3_tstrb,
    output [C_OUTPUT_BRAM_3_DMWIDTH-1:0] m_axis_bram_3_tdata,
    input m_axis_bram_3_tready,
    input [C_OUTPUT_BRAM_3_ADDR_WIDTH-1:0] ap_bram_oarg_3_addr0,
    input [C_OUTPUT_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_din0,
    output [C_OUTPUT_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_dout0,
    input ap_bram_oarg_3_clk0,
    input ap_bram_oarg_3_rst0,
    input [C_OUTPUT_BRAM_3_WIDTH/8-1:0] ap_bram_oarg_3_we0,
    input ap_bram_oarg_3_en0,
    input [C_OUTPUT_BRAM_3_ADDR_WIDTH-1:0] ap_bram_oarg_3_addr1,
    input [C_OUTPUT_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_din1,
    output [C_OUTPUT_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_dout1,
    input ap_bram_oarg_3_clk1,
    input ap_bram_oarg_3_rst1,
    input [C_OUTPUT_BRAM_3_WIDTH/8-1:0] ap_bram_oarg_3_we1,
    input ap_bram_oarg_3_en1,
    //out AXI-Stream output interface 4
    output m_axis_bram_4_tlast,
    output m_axis_bram_4_tvalid,
    output [C_OUTPUT_BRAM_4_DMWIDTH/8-1:0] m_axis_bram_4_tkeep,
    output [C_OUTPUT_BRAM_4_DMWIDTH/8-1:0] m_axis_bram_4_tstrb,
    output [C_OUTPUT_BRAM_4_DMWIDTH-1:0] m_axis_bram_4_tdata,
    input m_axis_bram_4_tready,
    input [C_OUTPUT_BRAM_4_ADDR_WIDTH-1:0] ap_bram_oarg_4_addr0,
    input [C_OUTPUT_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_din0,
    output [C_OUTPUT_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_dout0,
    input ap_bram_oarg_4_clk0,
    input ap_bram_oarg_4_rst0,
    input [C_OUTPUT_BRAM_4_WIDTH/8-1:0] ap_bram_oarg_4_we0,
    input ap_bram_oarg_4_en0,
    input [C_OUTPUT_BRAM_4_ADDR_WIDTH-1:0] ap_bram_oarg_4_addr1,
    input [C_OUTPUT_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_din1,
    output [C_OUTPUT_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_dout1,
    input ap_bram_oarg_4_clk1,
    input ap_bram_oarg_4_rst1,
    input [C_OUTPUT_BRAM_4_WIDTH/8-1:0] ap_bram_oarg_4_we1,
    input ap_bram_oarg_4_en1,
    //out AXI-Stream output interface 5
    output m_axis_bram_5_tlast,
    output m_axis_bram_5_tvalid,
    output [C_OUTPUT_BRAM_5_DMWIDTH/8-1:0] m_axis_bram_5_tkeep,
    output [C_OUTPUT_BRAM_5_DMWIDTH/8-1:0] m_axis_bram_5_tstrb,
    output [C_OUTPUT_BRAM_5_DMWIDTH-1:0] m_axis_bram_5_tdata,
    input m_axis_bram_5_tready,
    input [C_OUTPUT_BRAM_5_ADDR_WIDTH-1:0] ap_bram_oarg_5_addr0,
    input [C_OUTPUT_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_din0,
    output [C_OUTPUT_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_dout0,
    input ap_bram_oarg_5_clk0,
    input ap_bram_oarg_5_rst0,
    input [C_OUTPUT_BRAM_5_WIDTH/8-1:0] ap_bram_oarg_5_we0,
    input ap_bram_oarg_5_en0,
    input [C_OUTPUT_BRAM_5_ADDR_WIDTH-1:0] ap_bram_oarg_5_addr1,
    input [C_OUTPUT_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_din1,
    output [C_OUTPUT_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_dout1,
    input ap_bram_oarg_5_clk1,
    input ap_bram_oarg_5_rst1,
    input [C_OUTPUT_BRAM_5_WIDTH/8-1:0] ap_bram_oarg_5_we1,
    input ap_bram_oarg_5_en1,
    //out AXI-Stream output interface 6
    output m_axis_bram_6_tlast,
    output m_axis_bram_6_tvalid,
    output [C_OUTPUT_BRAM_6_DMWIDTH/8-1:0] m_axis_bram_6_tkeep,
    output [C_OUTPUT_BRAM_6_DMWIDTH/8-1:0] m_axis_bram_6_tstrb,
    output [C_OUTPUT_BRAM_6_DMWIDTH-1:0] m_axis_bram_6_tdata,
    input m_axis_bram_6_tready,
    input [C_OUTPUT_BRAM_6_ADDR_WIDTH-1:0] ap_bram_oarg_6_addr0,
    input [C_OUTPUT_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_din0,
    output [C_OUTPUT_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_dout0,
    input ap_bram_oarg_6_clk0,
    input ap_bram_oarg_6_rst0,
    input [C_OUTPUT_BRAM_6_WIDTH/8-1:0] ap_bram_oarg_6_we0,
    input ap_bram_oarg_6_en0,
    input [C_OUTPUT_BRAM_6_ADDR_WIDTH-1:0] ap_bram_oarg_6_addr1,
    input [C_OUTPUT_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_din1,
    output [C_OUTPUT_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_dout1,
    input ap_bram_oarg_6_clk1,
    input ap_bram_oarg_6_rst1,
    input [C_OUTPUT_BRAM_6_WIDTH/8-1:0] ap_bram_oarg_6_we1,
    input ap_bram_oarg_6_en1,
    //out AXI-Stream output interface 7
    output m_axis_bram_7_tlast,
    output m_axis_bram_7_tvalid,
    output [C_OUTPUT_BRAM_7_DMWIDTH/8-1:0] m_axis_bram_7_tkeep,
    output [C_OUTPUT_BRAM_7_DMWIDTH/8-1:0] m_axis_bram_7_tstrb,
    output [C_OUTPUT_BRAM_7_DMWIDTH-1:0] m_axis_bram_7_tdata,
    input m_axis_bram_7_tready,
    input [C_OUTPUT_BRAM_7_ADDR_WIDTH-1:0] ap_bram_oarg_7_addr0,
    input [C_OUTPUT_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_din0,
    output [C_OUTPUT_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_dout0,
    input ap_bram_oarg_7_clk0,
    input ap_bram_oarg_7_rst0,
    input [C_OUTPUT_BRAM_7_WIDTH/8-1:0] ap_bram_oarg_7_we0,
    input ap_bram_oarg_7_en0,
    input [C_OUTPUT_BRAM_7_ADDR_WIDTH-1:0] ap_bram_oarg_7_addr1,
    input [C_OUTPUT_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_din1,
    output [C_OUTPUT_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_dout1,
    input ap_bram_oarg_7_clk1,
    input ap_bram_oarg_7_rst1,
    input [C_OUTPUT_BRAM_7_WIDTH/8-1:0] ap_bram_oarg_7_we1,
    input ap_bram_oarg_7_en1,
    //out AXI-Stream output interface 8
    output m_axis_bram_8_tlast,
    output m_axis_bram_8_tvalid,
    output [C_OUTPUT_BRAM_8_DMWIDTH/8-1:0] m_axis_bram_8_tkeep,
    output [C_OUTPUT_BRAM_8_DMWIDTH/8-1:0] m_axis_bram_8_tstrb,
    output [C_OUTPUT_BRAM_8_DMWIDTH-1:0] m_axis_bram_8_tdata,
    input m_axis_bram_8_tready,
    input [C_OUTPUT_BRAM_8_ADDR_WIDTH-1:0] ap_bram_oarg_8_addr0,
    input [C_OUTPUT_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_din0,
    output [C_OUTPUT_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_dout0,
    input ap_bram_oarg_8_clk0,
    input ap_bram_oarg_8_rst0,
    input [C_OUTPUT_BRAM_8_WIDTH/8-1:0] ap_bram_oarg_8_we0,
    input ap_bram_oarg_8_en0,
    input [C_OUTPUT_BRAM_8_ADDR_WIDTH-1:0] ap_bram_oarg_8_addr1,
    input [C_OUTPUT_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_din1,
    output [C_OUTPUT_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_dout1,
    input ap_bram_oarg_8_clk1,
    input ap_bram_oarg_8_rst1,
    input [C_OUTPUT_BRAM_8_WIDTH/8-1:0] ap_bram_oarg_8_we1,
    input ap_bram_oarg_8_en1,
    //out AXI-Stream output interface 9
    output m_axis_bram_9_tlast,
    output m_axis_bram_9_tvalid,
    output [C_OUTPUT_BRAM_9_DMWIDTH/8-1:0] m_axis_bram_9_tkeep,
    output [C_OUTPUT_BRAM_9_DMWIDTH/8-1:0] m_axis_bram_9_tstrb,
    output [C_OUTPUT_BRAM_9_DMWIDTH-1:0] m_axis_bram_9_tdata,
    input m_axis_bram_9_tready,
    input [C_OUTPUT_BRAM_9_ADDR_WIDTH-1:0] ap_bram_oarg_9_addr0,
    input [C_OUTPUT_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_din0,
    output [C_OUTPUT_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_dout0,
    input ap_bram_oarg_9_clk0,
    input ap_bram_oarg_9_rst0,
    input [C_OUTPUT_BRAM_9_WIDTH/8-1:0] ap_bram_oarg_9_we0,
    input ap_bram_oarg_9_en0,
    input [C_OUTPUT_BRAM_9_ADDR_WIDTH-1:0] ap_bram_oarg_9_addr1,
    input [C_OUTPUT_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_din1,
    output [C_OUTPUT_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_dout1,
    input ap_bram_oarg_9_clk1,
    input ap_bram_oarg_9_rst1,
    input [C_OUTPUT_BRAM_9_WIDTH/8-1:0] ap_bram_oarg_9_we1,
    input ap_bram_oarg_9_en1,
    //out AXI-Stream output interface 10
    output m_axis_bram_10_tlast,
    output m_axis_bram_10_tvalid,
    output [C_OUTPUT_BRAM_10_DMWIDTH/8-1:0] m_axis_bram_10_tkeep,
    output [C_OUTPUT_BRAM_10_DMWIDTH/8-1:0] m_axis_bram_10_tstrb,
    output [C_OUTPUT_BRAM_10_DMWIDTH-1:0] m_axis_bram_10_tdata,
    input m_axis_bram_10_tready,
    input [C_OUTPUT_BRAM_10_ADDR_WIDTH-1:0] ap_bram_oarg_10_addr0,
    input [C_OUTPUT_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_din0,
    output [C_OUTPUT_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_dout0,
    input ap_bram_oarg_10_clk0,
    input ap_bram_oarg_10_rst0,
    input [C_OUTPUT_BRAM_10_WIDTH/8-1:0] ap_bram_oarg_10_we0,
    input ap_bram_oarg_10_en0,
    input [C_OUTPUT_BRAM_10_ADDR_WIDTH-1:0] ap_bram_oarg_10_addr1,
    input [C_OUTPUT_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_din1,
    output [C_OUTPUT_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_dout1,
    input ap_bram_oarg_10_clk1,
    input ap_bram_oarg_10_rst1,
    input [C_OUTPUT_BRAM_10_WIDTH/8-1:0] ap_bram_oarg_10_we1,
    input ap_bram_oarg_10_en1,
    //out AXI-Stream output interface 11
    output m_axis_bram_11_tlast,
    output m_axis_bram_11_tvalid,
    output [C_OUTPUT_BRAM_11_DMWIDTH/8-1:0] m_axis_bram_11_tkeep,
    output [C_OUTPUT_BRAM_11_DMWIDTH/8-1:0] m_axis_bram_11_tstrb,
    output [C_OUTPUT_BRAM_11_DMWIDTH-1:0] m_axis_bram_11_tdata,
    input m_axis_bram_11_tready,
    input [C_OUTPUT_BRAM_11_ADDR_WIDTH-1:0] ap_bram_oarg_11_addr0,
    input [C_OUTPUT_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_din0,
    output [C_OUTPUT_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_dout0,
    input ap_bram_oarg_11_clk0,
    input ap_bram_oarg_11_rst0,
    input [C_OUTPUT_BRAM_11_WIDTH/8-1:0] ap_bram_oarg_11_we0,
    input ap_bram_oarg_11_en0,
    input [C_OUTPUT_BRAM_11_ADDR_WIDTH-1:0] ap_bram_oarg_11_addr1,
    input [C_OUTPUT_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_din1,
    output [C_OUTPUT_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_dout1,
    input ap_bram_oarg_11_clk1,
    input ap_bram_oarg_11_rst1,
    input [C_OUTPUT_BRAM_11_WIDTH/8-1:0] ap_bram_oarg_11_we1,
    input ap_bram_oarg_11_en1,
    //out AXI-Stream output interface 12
    output m_axis_bram_12_tlast,
    output m_axis_bram_12_tvalid,
    output [C_OUTPUT_BRAM_12_DMWIDTH/8-1:0] m_axis_bram_12_tkeep,
    output [C_OUTPUT_BRAM_12_DMWIDTH/8-1:0] m_axis_bram_12_tstrb,
    output [C_OUTPUT_BRAM_12_DMWIDTH-1:0] m_axis_bram_12_tdata,
    input m_axis_bram_12_tready,
    input [C_OUTPUT_BRAM_12_ADDR_WIDTH-1:0] ap_bram_oarg_12_addr0,
    input [C_OUTPUT_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_din0,
    output [C_OUTPUT_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_dout0,
    input ap_bram_oarg_12_clk0,
    input ap_bram_oarg_12_rst0,
    input [C_OUTPUT_BRAM_12_WIDTH/8-1:0] ap_bram_oarg_12_we0,
    input ap_bram_oarg_12_en0,
    input [C_OUTPUT_BRAM_12_ADDR_WIDTH-1:0] ap_bram_oarg_12_addr1,
    input [C_OUTPUT_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_din1,
    output [C_OUTPUT_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_dout1,
    input ap_bram_oarg_12_clk1,
    input ap_bram_oarg_12_rst1,
    input [C_OUTPUT_BRAM_12_WIDTH/8-1:0] ap_bram_oarg_12_we1,
    input ap_bram_oarg_12_en1,
    //out AXI-Stream output interface 13
    output m_axis_bram_13_tlast,
    output m_axis_bram_13_tvalid,
    output [C_OUTPUT_BRAM_13_DMWIDTH/8-1:0] m_axis_bram_13_tkeep,
    output [C_OUTPUT_BRAM_13_DMWIDTH/8-1:0] m_axis_bram_13_tstrb,
    output [C_OUTPUT_BRAM_13_DMWIDTH-1:0] m_axis_bram_13_tdata,
    input m_axis_bram_13_tready,
    input [C_OUTPUT_BRAM_13_ADDR_WIDTH-1:0] ap_bram_oarg_13_addr0,
    input [C_OUTPUT_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_din0,
    output [C_OUTPUT_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_dout0,
    input ap_bram_oarg_13_clk0,
    input ap_bram_oarg_13_rst0,
    input [C_OUTPUT_BRAM_13_WIDTH/8-1:0] ap_bram_oarg_13_we0,
    input ap_bram_oarg_13_en0,
    input [C_OUTPUT_BRAM_13_ADDR_WIDTH-1:0] ap_bram_oarg_13_addr1,
    input [C_OUTPUT_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_din1,
    output [C_OUTPUT_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_dout1,
    input ap_bram_oarg_13_clk1,
    input ap_bram_oarg_13_rst1,
    input [C_OUTPUT_BRAM_13_WIDTH/8-1:0] ap_bram_oarg_13_we1,
    input ap_bram_oarg_13_en1,
    //out AXI-Stream output interface 14
    output m_axis_bram_14_tlast,
    output m_axis_bram_14_tvalid,
    output [C_OUTPUT_BRAM_14_DMWIDTH/8-1:0] m_axis_bram_14_tkeep,
    output [C_OUTPUT_BRAM_14_DMWIDTH/8-1:0] m_axis_bram_14_tstrb,
    output [C_OUTPUT_BRAM_14_DMWIDTH-1:0] m_axis_bram_14_tdata,
    input m_axis_bram_14_tready,
    input [C_OUTPUT_BRAM_14_ADDR_WIDTH-1:0] ap_bram_oarg_14_addr0,
    input [C_OUTPUT_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_din0,
    output [C_OUTPUT_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_dout0,
    input ap_bram_oarg_14_clk0,
    input ap_bram_oarg_14_rst0,
    input [C_OUTPUT_BRAM_14_WIDTH/8-1:0] ap_bram_oarg_14_we0,
    input ap_bram_oarg_14_en0,
    input [C_OUTPUT_BRAM_14_ADDR_WIDTH-1:0] ap_bram_oarg_14_addr1,
    input [C_OUTPUT_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_din1,
    output [C_OUTPUT_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_dout1,
    input ap_bram_oarg_14_clk1,
    input ap_bram_oarg_14_rst1,
    input [C_OUTPUT_BRAM_14_WIDTH/8-1:0] ap_bram_oarg_14_we1,
    input ap_bram_oarg_14_en1,
    //out AXI-Stream output interface 15
    output m_axis_bram_15_tlast,
    output m_axis_bram_15_tvalid,
    output [C_OUTPUT_BRAM_15_DMWIDTH/8-1:0] m_axis_bram_15_tkeep,
    output [C_OUTPUT_BRAM_15_DMWIDTH/8-1:0] m_axis_bram_15_tstrb,
    output [C_OUTPUT_BRAM_15_DMWIDTH-1:0] m_axis_bram_15_tdata,
    input m_axis_bram_15_tready,
    input [C_OUTPUT_BRAM_15_ADDR_WIDTH-1:0] ap_bram_oarg_15_addr0,
    input [C_OUTPUT_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_din0,
    output [C_OUTPUT_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_dout0,
    input ap_bram_oarg_15_clk0,
    input ap_bram_oarg_15_rst0,
    input [C_OUTPUT_BRAM_15_WIDTH/8-1:0] ap_bram_oarg_15_we0,
    input ap_bram_oarg_15_en0,
    input [C_OUTPUT_BRAM_15_ADDR_WIDTH-1:0] ap_bram_oarg_15_addr1,
    input [C_OUTPUT_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_din1,
    output [C_OUTPUT_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_dout1,
    input ap_bram_oarg_15_clk1,
    input ap_bram_oarg_15_rst1,
    input [C_OUTPUT_BRAM_15_WIDTH/8-1:0] ap_bram_oarg_15_we1,
    input ap_bram_oarg_15_en1,
    //out AXI-Stream output interface 16
    output m_axis_bram_16_tlast,
    output m_axis_bram_16_tvalid,
    output [C_OUTPUT_BRAM_16_DMWIDTH/8-1:0] m_axis_bram_16_tkeep,
    output [C_OUTPUT_BRAM_16_DMWIDTH/8-1:0] m_axis_bram_16_tstrb,
    output [C_OUTPUT_BRAM_16_DMWIDTH-1:0] m_axis_bram_16_tdata,
    input m_axis_bram_16_tready,
    input [C_OUTPUT_BRAM_16_ADDR_WIDTH-1:0] ap_bram_oarg_16_addr0,
    input [C_OUTPUT_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_din0,
    output [C_OUTPUT_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_dout0,
    input ap_bram_oarg_16_clk0,
    input ap_bram_oarg_16_rst0,
    input [C_OUTPUT_BRAM_16_WIDTH/8-1:0] ap_bram_oarg_16_we0,
    input ap_bram_oarg_16_en0,
    input [C_OUTPUT_BRAM_16_ADDR_WIDTH-1:0] ap_bram_oarg_16_addr1,
    input [C_OUTPUT_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_din1,
    output [C_OUTPUT_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_dout1,
    input ap_bram_oarg_16_clk1,
    input ap_bram_oarg_16_rst1,
    input [C_OUTPUT_BRAM_16_WIDTH/8-1:0] ap_bram_oarg_16_we1,
    input ap_bram_oarg_16_en1,
    //out AXI-Stream output interface 17
    output m_axis_bram_17_tlast,
    output m_axis_bram_17_tvalid,
    output [C_OUTPUT_BRAM_17_DMWIDTH/8-1:0] m_axis_bram_17_tkeep,
    output [C_OUTPUT_BRAM_17_DMWIDTH/8-1:0] m_axis_bram_17_tstrb,
    output [C_OUTPUT_BRAM_17_DMWIDTH-1:0] m_axis_bram_17_tdata,
    input m_axis_bram_17_tready,
    input [C_OUTPUT_BRAM_17_ADDR_WIDTH-1:0] ap_bram_oarg_17_addr0,
    input [C_OUTPUT_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_din0,
    output [C_OUTPUT_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_dout0,
    input ap_bram_oarg_17_clk0,
    input ap_bram_oarg_17_rst0,
    input [C_OUTPUT_BRAM_17_WIDTH/8-1:0] ap_bram_oarg_17_we0,
    input ap_bram_oarg_17_en0,
    input [C_OUTPUT_BRAM_17_ADDR_WIDTH-1:0] ap_bram_oarg_17_addr1,
    input [C_OUTPUT_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_din1,
    output [C_OUTPUT_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_dout1,
    input ap_bram_oarg_17_clk1,
    input ap_bram_oarg_17_rst1,
    input [C_OUTPUT_BRAM_17_WIDTH/8-1:0] ap_bram_oarg_17_we1,
    input ap_bram_oarg_17_en1,
    //out AXI-Stream output interface 18
    output m_axis_bram_18_tlast,
    output m_axis_bram_18_tvalid,
    output [C_OUTPUT_BRAM_18_DMWIDTH/8-1:0] m_axis_bram_18_tkeep,
    output [C_OUTPUT_BRAM_18_DMWIDTH/8-1:0] m_axis_bram_18_tstrb,
    output [C_OUTPUT_BRAM_18_DMWIDTH-1:0] m_axis_bram_18_tdata,
    input m_axis_bram_18_tready,
    input [C_OUTPUT_BRAM_18_ADDR_WIDTH-1:0] ap_bram_oarg_18_addr0,
    input [C_OUTPUT_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_din0,
    output [C_OUTPUT_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_dout0,
    input ap_bram_oarg_18_clk0,
    input ap_bram_oarg_18_rst0,
    input [C_OUTPUT_BRAM_18_WIDTH/8-1:0] ap_bram_oarg_18_we0,
    input ap_bram_oarg_18_en0,
    input [C_OUTPUT_BRAM_18_ADDR_WIDTH-1:0] ap_bram_oarg_18_addr1,
    input [C_OUTPUT_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_din1,
    output [C_OUTPUT_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_dout1,
    input ap_bram_oarg_18_clk1,
    input ap_bram_oarg_18_rst1,
    input [C_OUTPUT_BRAM_18_WIDTH/8-1:0] ap_bram_oarg_18_we1,
    input ap_bram_oarg_18_en1,
    //out AXI-Stream output interface 19
    output m_axis_bram_19_tlast,
    output m_axis_bram_19_tvalid,
    output [C_OUTPUT_BRAM_19_DMWIDTH/8-1:0] m_axis_bram_19_tkeep,
    output [C_OUTPUT_BRAM_19_DMWIDTH/8-1:0] m_axis_bram_19_tstrb,
    output [C_OUTPUT_BRAM_19_DMWIDTH-1:0] m_axis_bram_19_tdata,
    input m_axis_bram_19_tready,
    input [C_OUTPUT_BRAM_19_ADDR_WIDTH-1:0] ap_bram_oarg_19_addr0,
    input [C_OUTPUT_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_din0,
    output [C_OUTPUT_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_dout0,
    input ap_bram_oarg_19_clk0,
    input ap_bram_oarg_19_rst0,
    input [C_OUTPUT_BRAM_19_WIDTH/8-1:0] ap_bram_oarg_19_we0,
    input ap_bram_oarg_19_en0,
    input [C_OUTPUT_BRAM_19_ADDR_WIDTH-1:0] ap_bram_oarg_19_addr1,
    input [C_OUTPUT_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_din1,
    output [C_OUTPUT_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_dout1,
    input ap_bram_oarg_19_clk1,
    input ap_bram_oarg_19_rst1,
    input [C_OUTPUT_BRAM_19_WIDTH/8-1:0] ap_bram_oarg_19_we1,
    input ap_bram_oarg_19_en1,
    //out AXI-Stream output interface 20
    output m_axis_bram_20_tlast,
    output m_axis_bram_20_tvalid,
    output [C_OUTPUT_BRAM_20_DMWIDTH/8-1:0] m_axis_bram_20_tkeep,
    output [C_OUTPUT_BRAM_20_DMWIDTH/8-1:0] m_axis_bram_20_tstrb,
    output [C_OUTPUT_BRAM_20_DMWIDTH-1:0] m_axis_bram_20_tdata,
    input m_axis_bram_20_tready,
    input [C_OUTPUT_BRAM_20_ADDR_WIDTH-1:0] ap_bram_oarg_20_addr0,
    input [C_OUTPUT_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_din0,
    output [C_OUTPUT_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_dout0,
    input ap_bram_oarg_20_clk0,
    input ap_bram_oarg_20_rst0,
    input [C_OUTPUT_BRAM_20_WIDTH/8-1:0] ap_bram_oarg_20_we0,
    input ap_bram_oarg_20_en0,
    input [C_OUTPUT_BRAM_20_ADDR_WIDTH-1:0] ap_bram_oarg_20_addr1,
    input [C_OUTPUT_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_din1,
    output [C_OUTPUT_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_dout1,
    input ap_bram_oarg_20_clk1,
    input ap_bram_oarg_20_rst1,
    input [C_OUTPUT_BRAM_20_WIDTH/8-1:0] ap_bram_oarg_20_we1,
    input ap_bram_oarg_20_en1,
    //out AXI-Stream output interface 21
    output m_axis_bram_21_tlast,
    output m_axis_bram_21_tvalid,
    output [C_OUTPUT_BRAM_21_DMWIDTH/8-1:0] m_axis_bram_21_tkeep,
    output [C_OUTPUT_BRAM_21_DMWIDTH/8-1:0] m_axis_bram_21_tstrb,
    output [C_OUTPUT_BRAM_21_DMWIDTH-1:0] m_axis_bram_21_tdata,
    input m_axis_bram_21_tready,
    input [C_OUTPUT_BRAM_21_ADDR_WIDTH-1:0] ap_bram_oarg_21_addr0,
    input [C_OUTPUT_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_din0,
    output [C_OUTPUT_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_dout0,
    input ap_bram_oarg_21_clk0,
    input ap_bram_oarg_21_rst0,
    input [C_OUTPUT_BRAM_21_WIDTH/8-1:0] ap_bram_oarg_21_we0,
    input ap_bram_oarg_21_en0,
    input [C_OUTPUT_BRAM_21_ADDR_WIDTH-1:0] ap_bram_oarg_21_addr1,
    input [C_OUTPUT_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_din1,
    output [C_OUTPUT_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_dout1,
    input ap_bram_oarg_21_clk1,
    input ap_bram_oarg_21_rst1,
    input [C_OUTPUT_BRAM_21_WIDTH/8-1:0] ap_bram_oarg_21_we1,
    input ap_bram_oarg_21_en1,
    //out AXI-Stream output interface 22
    output m_axis_bram_22_tlast,
    output m_axis_bram_22_tvalid,
    output [C_OUTPUT_BRAM_22_DMWIDTH/8-1:0] m_axis_bram_22_tkeep,
    output [C_OUTPUT_BRAM_22_DMWIDTH/8-1:0] m_axis_bram_22_tstrb,
    output [C_OUTPUT_BRAM_22_DMWIDTH-1:0] m_axis_bram_22_tdata,
    input m_axis_bram_22_tready,
    input [C_OUTPUT_BRAM_22_ADDR_WIDTH-1:0] ap_bram_oarg_22_addr0,
    input [C_OUTPUT_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_din0,
    output [C_OUTPUT_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_dout0,
    input ap_bram_oarg_22_clk0,
    input ap_bram_oarg_22_rst0,
    input [C_OUTPUT_BRAM_22_WIDTH/8-1:0] ap_bram_oarg_22_we0,
    input ap_bram_oarg_22_en0,
    input [C_OUTPUT_BRAM_22_ADDR_WIDTH-1:0] ap_bram_oarg_22_addr1,
    input [C_OUTPUT_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_din1,
    output [C_OUTPUT_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_dout1,
    input ap_bram_oarg_22_clk1,
    input ap_bram_oarg_22_rst1,
    input [C_OUTPUT_BRAM_22_WIDTH/8-1:0] ap_bram_oarg_22_we1,
    input ap_bram_oarg_22_en1,
    //out AXI-Stream output interface 23
    output m_axis_bram_23_tlast,
    output m_axis_bram_23_tvalid,
    output [C_OUTPUT_BRAM_23_DMWIDTH/8-1:0] m_axis_bram_23_tkeep,
    output [C_OUTPUT_BRAM_23_DMWIDTH/8-1:0] m_axis_bram_23_tstrb,
    output [C_OUTPUT_BRAM_23_DMWIDTH-1:0] m_axis_bram_23_tdata,
    input m_axis_bram_23_tready,
    input [C_OUTPUT_BRAM_23_ADDR_WIDTH-1:0] ap_bram_oarg_23_addr0,
    input [C_OUTPUT_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_din0,
    output [C_OUTPUT_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_dout0,
    input ap_bram_oarg_23_clk0,
    input ap_bram_oarg_23_rst0,
    input [C_OUTPUT_BRAM_23_WIDTH/8-1:0] ap_bram_oarg_23_we0,
    input ap_bram_oarg_23_en0,
    input [C_OUTPUT_BRAM_23_ADDR_WIDTH-1:0] ap_bram_oarg_23_addr1,
    input [C_OUTPUT_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_din1,
    output [C_OUTPUT_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_dout1,
    input ap_bram_oarg_23_clk1,
    input ap_bram_oarg_23_rst1,
    input [C_OUTPUT_BRAM_23_WIDTH/8-1:0] ap_bram_oarg_23_we1,
    input ap_bram_oarg_23_en1,
    //out AXI-Stream output interface 24
    output m_axis_bram_24_tlast,
    output m_axis_bram_24_tvalid,
    output [C_OUTPUT_BRAM_24_DMWIDTH/8-1:0] m_axis_bram_24_tkeep,
    output [C_OUTPUT_BRAM_24_DMWIDTH/8-1:0] m_axis_bram_24_tstrb,
    output [C_OUTPUT_BRAM_24_DMWIDTH-1:0] m_axis_bram_24_tdata,
    input m_axis_bram_24_tready,
    input [C_OUTPUT_BRAM_24_ADDR_WIDTH-1:0] ap_bram_oarg_24_addr0,
    input [C_OUTPUT_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_din0,
    output [C_OUTPUT_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_dout0,
    input ap_bram_oarg_24_clk0,
    input ap_bram_oarg_24_rst0,
    input [C_OUTPUT_BRAM_24_WIDTH/8-1:0] ap_bram_oarg_24_we0,
    input ap_bram_oarg_24_en0,
    input [C_OUTPUT_BRAM_24_ADDR_WIDTH-1:0] ap_bram_oarg_24_addr1,
    input [C_OUTPUT_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_din1,
    output [C_OUTPUT_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_dout1,
    input ap_bram_oarg_24_clk1,
    input ap_bram_oarg_24_rst1,
    input [C_OUTPUT_BRAM_24_WIDTH/8-1:0] ap_bram_oarg_24_we1,
    input ap_bram_oarg_24_en1,
    //out AXI-Stream output interface 25
    output m_axis_bram_25_tlast,
    output m_axis_bram_25_tvalid,
    output [C_OUTPUT_BRAM_25_DMWIDTH/8-1:0] m_axis_bram_25_tkeep,
    output [C_OUTPUT_BRAM_25_DMWIDTH/8-1:0] m_axis_bram_25_tstrb,
    output [C_OUTPUT_BRAM_25_DMWIDTH-1:0] m_axis_bram_25_tdata,
    input m_axis_bram_25_tready,
    input [C_OUTPUT_BRAM_25_ADDR_WIDTH-1:0] ap_bram_oarg_25_addr0,
    input [C_OUTPUT_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_din0,
    output [C_OUTPUT_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_dout0,
    input ap_bram_oarg_25_clk0,
    input ap_bram_oarg_25_rst0,
    input [C_OUTPUT_BRAM_25_WIDTH/8-1:0] ap_bram_oarg_25_we0,
    input ap_bram_oarg_25_en0,
    input [C_OUTPUT_BRAM_25_ADDR_WIDTH-1:0] ap_bram_oarg_25_addr1,
    input [C_OUTPUT_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_din1,
    output [C_OUTPUT_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_dout1,
    input ap_bram_oarg_25_clk1,
    input ap_bram_oarg_25_rst1,
    input [C_OUTPUT_BRAM_25_WIDTH/8-1:0] ap_bram_oarg_25_we1,
    input ap_bram_oarg_25_en1,
    //out AXI-Stream output interface 26
    output m_axis_bram_26_tlast,
    output m_axis_bram_26_tvalid,
    output [C_OUTPUT_BRAM_26_DMWIDTH/8-1:0] m_axis_bram_26_tkeep,
    output [C_OUTPUT_BRAM_26_DMWIDTH/8-1:0] m_axis_bram_26_tstrb,
    output [C_OUTPUT_BRAM_26_DMWIDTH-1:0] m_axis_bram_26_tdata,
    input m_axis_bram_26_tready,
    input [C_OUTPUT_BRAM_26_ADDR_WIDTH-1:0] ap_bram_oarg_26_addr0,
    input [C_OUTPUT_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_din0,
    output [C_OUTPUT_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_dout0,
    input ap_bram_oarg_26_clk0,
    input ap_bram_oarg_26_rst0,
    input [C_OUTPUT_BRAM_26_WIDTH/8-1:0] ap_bram_oarg_26_we0,
    input ap_bram_oarg_26_en0,
    input [C_OUTPUT_BRAM_26_ADDR_WIDTH-1:0] ap_bram_oarg_26_addr1,
    input [C_OUTPUT_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_din1,
    output [C_OUTPUT_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_dout1,
    input ap_bram_oarg_26_clk1,
    input ap_bram_oarg_26_rst1,
    input [C_OUTPUT_BRAM_26_WIDTH/8-1:0] ap_bram_oarg_26_we1,
    input ap_bram_oarg_26_en1,
    //out AXI-Stream output interface 27
    output m_axis_bram_27_tlast,
    output m_axis_bram_27_tvalid,
    output [C_OUTPUT_BRAM_27_DMWIDTH/8-1:0] m_axis_bram_27_tkeep,
    output [C_OUTPUT_BRAM_27_DMWIDTH/8-1:0] m_axis_bram_27_tstrb,
    output [C_OUTPUT_BRAM_27_DMWIDTH-1:0] m_axis_bram_27_tdata,
    input m_axis_bram_27_tready,
    input [C_OUTPUT_BRAM_27_ADDR_WIDTH-1:0] ap_bram_oarg_27_addr0,
    input [C_OUTPUT_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_din0,
    output [C_OUTPUT_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_dout0,
    input ap_bram_oarg_27_clk0,
    input ap_bram_oarg_27_rst0,
    input [C_OUTPUT_BRAM_27_WIDTH/8-1:0] ap_bram_oarg_27_we0,
    input ap_bram_oarg_27_en0,
    input [C_OUTPUT_BRAM_27_ADDR_WIDTH-1:0] ap_bram_oarg_27_addr1,
    input [C_OUTPUT_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_din1,
    output [C_OUTPUT_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_dout1,
    input ap_bram_oarg_27_clk1,
    input ap_bram_oarg_27_rst1,
    input [C_OUTPUT_BRAM_27_WIDTH/8-1:0] ap_bram_oarg_27_we1,
    input ap_bram_oarg_27_en1,
    //out AXI-Stream output interface 28
    output m_axis_bram_28_tlast,
    output m_axis_bram_28_tvalid,
    output [C_OUTPUT_BRAM_28_DMWIDTH/8-1:0] m_axis_bram_28_tkeep,
    output [C_OUTPUT_BRAM_28_DMWIDTH/8-1:0] m_axis_bram_28_tstrb,
    output [C_OUTPUT_BRAM_28_DMWIDTH-1:0] m_axis_bram_28_tdata,
    input m_axis_bram_28_tready,
    input [C_OUTPUT_BRAM_28_ADDR_WIDTH-1:0] ap_bram_oarg_28_addr0,
    input [C_OUTPUT_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_din0,
    output [C_OUTPUT_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_dout0,
    input ap_bram_oarg_28_clk0,
    input ap_bram_oarg_28_rst0,
    input [C_OUTPUT_BRAM_28_WIDTH/8-1:0] ap_bram_oarg_28_we0,
    input ap_bram_oarg_28_en0,
    input [C_OUTPUT_BRAM_28_ADDR_WIDTH-1:0] ap_bram_oarg_28_addr1,
    input [C_OUTPUT_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_din1,
    output [C_OUTPUT_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_dout1,
    input ap_bram_oarg_28_clk1,
    input ap_bram_oarg_28_rst1,
    input [C_OUTPUT_BRAM_28_WIDTH/8-1:0] ap_bram_oarg_28_we1,
    input ap_bram_oarg_28_en1,
    //out AXI-Stream output interface 29
    output m_axis_bram_29_tlast,
    output m_axis_bram_29_tvalid,
    output [C_OUTPUT_BRAM_29_DMWIDTH/8-1:0] m_axis_bram_29_tkeep,
    output [C_OUTPUT_BRAM_29_DMWIDTH/8-1:0] m_axis_bram_29_tstrb,
    output [C_OUTPUT_BRAM_29_DMWIDTH-1:0] m_axis_bram_29_tdata,
    input m_axis_bram_29_tready,
    input [C_OUTPUT_BRAM_29_ADDR_WIDTH-1:0] ap_bram_oarg_29_addr0,
    input [C_OUTPUT_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_din0,
    output [C_OUTPUT_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_dout0,
    input ap_bram_oarg_29_clk0,
    input ap_bram_oarg_29_rst0,
    input [C_OUTPUT_BRAM_29_WIDTH/8-1:0] ap_bram_oarg_29_we0,
    input ap_bram_oarg_29_en0,
    input [C_OUTPUT_BRAM_29_ADDR_WIDTH-1:0] ap_bram_oarg_29_addr1,
    input [C_OUTPUT_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_din1,
    output [C_OUTPUT_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_dout1,
    input ap_bram_oarg_29_clk1,
    input ap_bram_oarg_29_rst1,
    input [C_OUTPUT_BRAM_29_WIDTH/8-1:0] ap_bram_oarg_29_we1,
    input ap_bram_oarg_29_en1,
    //out AXI-Stream output interface 30
    output m_axis_bram_30_tlast,
    output m_axis_bram_30_tvalid,
    output [C_OUTPUT_BRAM_30_DMWIDTH/8-1:0] m_axis_bram_30_tkeep,
    output [C_OUTPUT_BRAM_30_DMWIDTH/8-1:0] m_axis_bram_30_tstrb,
    output [C_OUTPUT_BRAM_30_DMWIDTH-1:0] m_axis_bram_30_tdata,
    input m_axis_bram_30_tready,
    input [C_OUTPUT_BRAM_30_ADDR_WIDTH-1:0] ap_bram_oarg_30_addr0,
    input [C_OUTPUT_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_din0,
    output [C_OUTPUT_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_dout0,
    input ap_bram_oarg_30_clk0,
    input ap_bram_oarg_30_rst0,
    input [C_OUTPUT_BRAM_30_WIDTH/8-1:0] ap_bram_oarg_30_we0,
    input ap_bram_oarg_30_en0,
    input [C_OUTPUT_BRAM_30_ADDR_WIDTH-1:0] ap_bram_oarg_30_addr1,
    input [C_OUTPUT_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_din1,
    output [C_OUTPUT_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_dout1,
    input ap_bram_oarg_30_clk1,
    input ap_bram_oarg_30_rst1,
    input [C_OUTPUT_BRAM_30_WIDTH/8-1:0] ap_bram_oarg_30_we1,
    input ap_bram_oarg_30_en1,
    //out AXI-Stream output interface 31
    output m_axis_bram_31_tlast,
    output m_axis_bram_31_tvalid,
    output [C_OUTPUT_BRAM_31_DMWIDTH/8-1:0] m_axis_bram_31_tkeep,
    output [C_OUTPUT_BRAM_31_DMWIDTH/8-1:0] m_axis_bram_31_tstrb,
    output [C_OUTPUT_BRAM_31_DMWIDTH-1:0] m_axis_bram_31_tdata,
    input m_axis_bram_31_tready,
    input [C_OUTPUT_BRAM_31_ADDR_WIDTH-1:0] ap_bram_oarg_31_addr0,
    input [C_OUTPUT_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_din0,
    output [C_OUTPUT_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_dout0,
    input ap_bram_oarg_31_clk0,
    input ap_bram_oarg_31_rst0,
    input [C_OUTPUT_BRAM_31_WIDTH/8-1:0] ap_bram_oarg_31_we0,
    input ap_bram_oarg_31_en0,
    input [C_OUTPUT_BRAM_31_ADDR_WIDTH-1:0] ap_bram_oarg_31_addr1,
    input [C_OUTPUT_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_din1,
    output [C_OUTPUT_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_dout1,
    input ap_bram_oarg_31_clk1,
    input ap_bram_oarg_31_rst1,
    input [C_OUTPUT_BRAM_31_WIDTH/8-1:0] ap_bram_oarg_31_we1,
    input ap_bram_oarg_31_en1,
    //out AXI-Stream output interface 32
    output m_axis_bram_32_tlast,
    output m_axis_bram_32_tvalid,
    output [C_OUTPUT_BRAM_32_DMWIDTH/8-1:0] m_axis_bram_32_tkeep,
    output [C_OUTPUT_BRAM_32_DMWIDTH/8-1:0] m_axis_bram_32_tstrb,
    output [C_OUTPUT_BRAM_32_DMWIDTH-1:0] m_axis_bram_32_tdata,
    input m_axis_bram_32_tready,
    input [C_OUTPUT_BRAM_32_ADDR_WIDTH-1:0] ap_bram_oarg_32_addr0,
    input [C_OUTPUT_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_din0,
    output [C_OUTPUT_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_dout0,
    input ap_bram_oarg_32_clk0,
    input ap_bram_oarg_32_rst0,
    input [C_OUTPUT_BRAM_32_WIDTH/8-1:0] ap_bram_oarg_32_we0,
    input ap_bram_oarg_32_en0,
    input [C_OUTPUT_BRAM_32_ADDR_WIDTH-1:0] ap_bram_oarg_32_addr1,
    input [C_OUTPUT_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_din1,
    output [C_OUTPUT_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_dout1,
    input ap_bram_oarg_32_clk1,
    input ap_bram_oarg_32_rst1,
    input [C_OUTPUT_BRAM_32_WIDTH/8-1:0] ap_bram_oarg_32_we1,
    input ap_bram_oarg_32_en1,
    //out AXI-Stream output interface 33
    output m_axis_bram_33_tlast,
    output m_axis_bram_33_tvalid,
    output [C_OUTPUT_BRAM_33_DMWIDTH/8-1:0] m_axis_bram_33_tkeep,
    output [C_OUTPUT_BRAM_33_DMWIDTH/8-1:0] m_axis_bram_33_tstrb,
    output [C_OUTPUT_BRAM_33_DMWIDTH-1:0] m_axis_bram_33_tdata,
    input m_axis_bram_33_tready,
    input [C_OUTPUT_BRAM_33_ADDR_WIDTH-1:0] ap_bram_oarg_33_addr0,
    input [C_OUTPUT_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_din0,
    output [C_OUTPUT_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_dout0,
    input ap_bram_oarg_33_clk0,
    input ap_bram_oarg_33_rst0,
    input [C_OUTPUT_BRAM_33_WIDTH/8-1:0] ap_bram_oarg_33_we0,
    input ap_bram_oarg_33_en0,
    input [C_OUTPUT_BRAM_33_ADDR_WIDTH-1:0] ap_bram_oarg_33_addr1,
    input [C_OUTPUT_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_din1,
    output [C_OUTPUT_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_dout1,
    input ap_bram_oarg_33_clk1,
    input ap_bram_oarg_33_rst1,
    input [C_OUTPUT_BRAM_33_WIDTH/8-1:0] ap_bram_oarg_33_we1,
    input ap_bram_oarg_33_en1,
    //out AXI-Stream output interface 34
    output m_axis_bram_34_tlast,
    output m_axis_bram_34_tvalid,
    output [C_OUTPUT_BRAM_34_DMWIDTH/8-1:0] m_axis_bram_34_tkeep,
    output [C_OUTPUT_BRAM_34_DMWIDTH/8-1:0] m_axis_bram_34_tstrb,
    output [C_OUTPUT_BRAM_34_DMWIDTH-1:0] m_axis_bram_34_tdata,
    input m_axis_bram_34_tready,
    input [C_OUTPUT_BRAM_34_ADDR_WIDTH-1:0] ap_bram_oarg_34_addr0,
    input [C_OUTPUT_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_din0,
    output [C_OUTPUT_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_dout0,
    input ap_bram_oarg_34_clk0,
    input ap_bram_oarg_34_rst0,
    input [C_OUTPUT_BRAM_34_WIDTH/8-1:0] ap_bram_oarg_34_we0,
    input ap_bram_oarg_34_en0,
    input [C_OUTPUT_BRAM_34_ADDR_WIDTH-1:0] ap_bram_oarg_34_addr1,
    input [C_OUTPUT_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_din1,
    output [C_OUTPUT_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_dout1,
    input ap_bram_oarg_34_clk1,
    input ap_bram_oarg_34_rst1,
    input [C_OUTPUT_BRAM_34_WIDTH/8-1:0] ap_bram_oarg_34_we1,
    input ap_bram_oarg_34_en1,
    //out AXI-Stream output interface 35
    output m_axis_bram_35_tlast,
    output m_axis_bram_35_tvalid,
    output [C_OUTPUT_BRAM_35_DMWIDTH/8-1:0] m_axis_bram_35_tkeep,
    output [C_OUTPUT_BRAM_35_DMWIDTH/8-1:0] m_axis_bram_35_tstrb,
    output [C_OUTPUT_BRAM_35_DMWIDTH-1:0] m_axis_bram_35_tdata,
    input m_axis_bram_35_tready,
    input [C_OUTPUT_BRAM_35_ADDR_WIDTH-1:0] ap_bram_oarg_35_addr0,
    input [C_OUTPUT_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_din0,
    output [C_OUTPUT_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_dout0,
    input ap_bram_oarg_35_clk0,
    input ap_bram_oarg_35_rst0,
    input [C_OUTPUT_BRAM_35_WIDTH/8-1:0] ap_bram_oarg_35_we0,
    input ap_bram_oarg_35_en0,
    input [C_OUTPUT_BRAM_35_ADDR_WIDTH-1:0] ap_bram_oarg_35_addr1,
    input [C_OUTPUT_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_din1,
    output [C_OUTPUT_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_dout1,
    input ap_bram_oarg_35_clk1,
    input ap_bram_oarg_35_rst1,
    input [C_OUTPUT_BRAM_35_WIDTH/8-1:0] ap_bram_oarg_35_we1,
    input ap_bram_oarg_35_en1,
    //out AXI-Stream output interface 36
    output m_axis_bram_36_tlast,
    output m_axis_bram_36_tvalid,
    output [C_OUTPUT_BRAM_36_DMWIDTH/8-1:0] m_axis_bram_36_tkeep,
    output [C_OUTPUT_BRAM_36_DMWIDTH/8-1:0] m_axis_bram_36_tstrb,
    output [C_OUTPUT_BRAM_36_DMWIDTH-1:0] m_axis_bram_36_tdata,
    input m_axis_bram_36_tready,
    input [C_OUTPUT_BRAM_36_ADDR_WIDTH-1:0] ap_bram_oarg_36_addr0,
    input [C_OUTPUT_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_din0,
    output [C_OUTPUT_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_dout0,
    input ap_bram_oarg_36_clk0,
    input ap_bram_oarg_36_rst0,
    input [C_OUTPUT_BRAM_36_WIDTH/8-1:0] ap_bram_oarg_36_we0,
    input ap_bram_oarg_36_en0,
    input [C_OUTPUT_BRAM_36_ADDR_WIDTH-1:0] ap_bram_oarg_36_addr1,
    input [C_OUTPUT_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_din1,
    output [C_OUTPUT_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_dout1,
    input ap_bram_oarg_36_clk1,
    input ap_bram_oarg_36_rst1,
    input [C_OUTPUT_BRAM_36_WIDTH/8-1:0] ap_bram_oarg_36_we1,
    input ap_bram_oarg_36_en1,
    //out AXI-Stream output interface 37
    output m_axis_bram_37_tlast,
    output m_axis_bram_37_tvalid,
    output [C_OUTPUT_BRAM_37_DMWIDTH/8-1:0] m_axis_bram_37_tkeep,
    output [C_OUTPUT_BRAM_37_DMWIDTH/8-1:0] m_axis_bram_37_tstrb,
    output [C_OUTPUT_BRAM_37_DMWIDTH-1:0] m_axis_bram_37_tdata,
    input m_axis_bram_37_tready,
    input [C_OUTPUT_BRAM_37_ADDR_WIDTH-1:0] ap_bram_oarg_37_addr0,
    input [C_OUTPUT_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_din0,
    output [C_OUTPUT_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_dout0,
    input ap_bram_oarg_37_clk0,
    input ap_bram_oarg_37_rst0,
    input [C_OUTPUT_BRAM_37_WIDTH/8-1:0] ap_bram_oarg_37_we0,
    input ap_bram_oarg_37_en0,
    input [C_OUTPUT_BRAM_37_ADDR_WIDTH-1:0] ap_bram_oarg_37_addr1,
    input [C_OUTPUT_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_din1,
    output [C_OUTPUT_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_dout1,
    input ap_bram_oarg_37_clk1,
    input ap_bram_oarg_37_rst1,
    input [C_OUTPUT_BRAM_37_WIDTH/8-1:0] ap_bram_oarg_37_we1,
    input ap_bram_oarg_37_en1,
    //out AXI-Stream output interface 38
    output m_axis_bram_38_tlast,
    output m_axis_bram_38_tvalid,
    output [C_OUTPUT_BRAM_38_DMWIDTH/8-1:0] m_axis_bram_38_tkeep,
    output [C_OUTPUT_BRAM_38_DMWIDTH/8-1:0] m_axis_bram_38_tstrb,
    output [C_OUTPUT_BRAM_38_DMWIDTH-1:0] m_axis_bram_38_tdata,
    input m_axis_bram_38_tready,
    input [C_OUTPUT_BRAM_38_ADDR_WIDTH-1:0] ap_bram_oarg_38_addr0,
    input [C_OUTPUT_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_din0,
    output [C_OUTPUT_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_dout0,
    input ap_bram_oarg_38_clk0,
    input ap_bram_oarg_38_rst0,
    input [C_OUTPUT_BRAM_38_WIDTH/8-1:0] ap_bram_oarg_38_we0,
    input ap_bram_oarg_38_en0,
    input [C_OUTPUT_BRAM_38_ADDR_WIDTH-1:0] ap_bram_oarg_38_addr1,
    input [C_OUTPUT_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_din1,
    output [C_OUTPUT_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_dout1,
    input ap_bram_oarg_38_clk1,
    input ap_bram_oarg_38_rst1,
    input [C_OUTPUT_BRAM_38_WIDTH/8-1:0] ap_bram_oarg_38_we1,
    input ap_bram_oarg_38_en1,
    //out AXI-Stream output interface 39
    output m_axis_bram_39_tlast,
    output m_axis_bram_39_tvalid,
    output [C_OUTPUT_BRAM_39_DMWIDTH/8-1:0] m_axis_bram_39_tkeep,
    output [C_OUTPUT_BRAM_39_DMWIDTH/8-1:0] m_axis_bram_39_tstrb,
    output [C_OUTPUT_BRAM_39_DMWIDTH-1:0] m_axis_bram_39_tdata,
    input m_axis_bram_39_tready,
    input [C_OUTPUT_BRAM_39_ADDR_WIDTH-1:0] ap_bram_oarg_39_addr0,
    input [C_OUTPUT_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_din0,
    output [C_OUTPUT_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_dout0,
    input ap_bram_oarg_39_clk0,
    input ap_bram_oarg_39_rst0,
    input [C_OUTPUT_BRAM_39_WIDTH/8-1:0] ap_bram_oarg_39_we0,
    input ap_bram_oarg_39_en0,
    input [C_OUTPUT_BRAM_39_ADDR_WIDTH-1:0] ap_bram_oarg_39_addr1,
    input [C_OUTPUT_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_din1,
    output [C_OUTPUT_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_dout1,
    input ap_bram_oarg_39_clk1,
    input ap_bram_oarg_39_rst1,
    input [C_OUTPUT_BRAM_39_WIDTH/8-1:0] ap_bram_oarg_39_we1,
    input ap_bram_oarg_39_en1,
    //out AXI-Stream output interface 40
    output m_axis_bram_40_tlast,
    output m_axis_bram_40_tvalid,
    output [C_OUTPUT_BRAM_40_DMWIDTH/8-1:0] m_axis_bram_40_tkeep,
    output [C_OUTPUT_BRAM_40_DMWIDTH/8-1:0] m_axis_bram_40_tstrb,
    output [C_OUTPUT_BRAM_40_DMWIDTH-1:0] m_axis_bram_40_tdata,
    input m_axis_bram_40_tready,
    input [C_OUTPUT_BRAM_40_ADDR_WIDTH-1:0] ap_bram_oarg_40_addr0,
    input [C_OUTPUT_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_din0,
    output [C_OUTPUT_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_dout0,
    input ap_bram_oarg_40_clk0,
    input ap_bram_oarg_40_rst0,
    input [C_OUTPUT_BRAM_40_WIDTH/8-1:0] ap_bram_oarg_40_we0,
    input ap_bram_oarg_40_en0,
    input [C_OUTPUT_BRAM_40_ADDR_WIDTH-1:0] ap_bram_oarg_40_addr1,
    input [C_OUTPUT_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_din1,
    output [C_OUTPUT_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_dout1,
    input ap_bram_oarg_40_clk1,
    input ap_bram_oarg_40_rst1,
    input [C_OUTPUT_BRAM_40_WIDTH/8-1:0] ap_bram_oarg_40_we1,
    input ap_bram_oarg_40_en1,
    //out AXI-Stream output interface 41
    output m_axis_bram_41_tlast,
    output m_axis_bram_41_tvalid,
    output [C_OUTPUT_BRAM_41_DMWIDTH/8-1:0] m_axis_bram_41_tkeep,
    output [C_OUTPUT_BRAM_41_DMWIDTH/8-1:0] m_axis_bram_41_tstrb,
    output [C_OUTPUT_BRAM_41_DMWIDTH-1:0] m_axis_bram_41_tdata,
    input m_axis_bram_41_tready,
    input [C_OUTPUT_BRAM_41_ADDR_WIDTH-1:0] ap_bram_oarg_41_addr0,
    input [C_OUTPUT_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_din0,
    output [C_OUTPUT_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_dout0,
    input ap_bram_oarg_41_clk0,
    input ap_bram_oarg_41_rst0,
    input [C_OUTPUT_BRAM_41_WIDTH/8-1:0] ap_bram_oarg_41_we0,
    input ap_bram_oarg_41_en0,
    input [C_OUTPUT_BRAM_41_ADDR_WIDTH-1:0] ap_bram_oarg_41_addr1,
    input [C_OUTPUT_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_din1,
    output [C_OUTPUT_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_dout1,
    input ap_bram_oarg_41_clk1,
    input ap_bram_oarg_41_rst1,
    input [C_OUTPUT_BRAM_41_WIDTH/8-1:0] ap_bram_oarg_41_we1,
    input ap_bram_oarg_41_en1,
    //out AXI-Stream output interface 42
    output m_axis_bram_42_tlast,
    output m_axis_bram_42_tvalid,
    output [C_OUTPUT_BRAM_42_DMWIDTH/8-1:0] m_axis_bram_42_tkeep,
    output [C_OUTPUT_BRAM_42_DMWIDTH/8-1:0] m_axis_bram_42_tstrb,
    output [C_OUTPUT_BRAM_42_DMWIDTH-1:0] m_axis_bram_42_tdata,
    input m_axis_bram_42_tready,
    input [C_OUTPUT_BRAM_42_ADDR_WIDTH-1:0] ap_bram_oarg_42_addr0,
    input [C_OUTPUT_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_din0,
    output [C_OUTPUT_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_dout0,
    input ap_bram_oarg_42_clk0,
    input ap_bram_oarg_42_rst0,
    input [C_OUTPUT_BRAM_42_WIDTH/8-1:0] ap_bram_oarg_42_we0,
    input ap_bram_oarg_42_en0,
    input [C_OUTPUT_BRAM_42_ADDR_WIDTH-1:0] ap_bram_oarg_42_addr1,
    input [C_OUTPUT_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_din1,
    output [C_OUTPUT_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_dout1,
    input ap_bram_oarg_42_clk1,
    input ap_bram_oarg_42_rst1,
    input [C_OUTPUT_BRAM_42_WIDTH/8-1:0] ap_bram_oarg_42_we1,
    input ap_bram_oarg_42_en1,
    //out AXI-Stream output interface 43
    output m_axis_bram_43_tlast,
    output m_axis_bram_43_tvalid,
    output [C_OUTPUT_BRAM_43_DMWIDTH/8-1:0] m_axis_bram_43_tkeep,
    output [C_OUTPUT_BRAM_43_DMWIDTH/8-1:0] m_axis_bram_43_tstrb,
    output [C_OUTPUT_BRAM_43_DMWIDTH-1:0] m_axis_bram_43_tdata,
    input m_axis_bram_43_tready,
    input [C_OUTPUT_BRAM_43_ADDR_WIDTH-1:0] ap_bram_oarg_43_addr0,
    input [C_OUTPUT_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_din0,
    output [C_OUTPUT_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_dout0,
    input ap_bram_oarg_43_clk0,
    input ap_bram_oarg_43_rst0,
    input [C_OUTPUT_BRAM_43_WIDTH/8-1:0] ap_bram_oarg_43_we0,
    input ap_bram_oarg_43_en0,
    input [C_OUTPUT_BRAM_43_ADDR_WIDTH-1:0] ap_bram_oarg_43_addr1,
    input [C_OUTPUT_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_din1,
    output [C_OUTPUT_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_dout1,
    input ap_bram_oarg_43_clk1,
    input ap_bram_oarg_43_rst1,
    input [C_OUTPUT_BRAM_43_WIDTH/8-1:0] ap_bram_oarg_43_we1,
    input ap_bram_oarg_43_en1,
    //out AXI-Stream output interface 44
    output m_axis_bram_44_tlast,
    output m_axis_bram_44_tvalid,
    output [C_OUTPUT_BRAM_44_DMWIDTH/8-1:0] m_axis_bram_44_tkeep,
    output [C_OUTPUT_BRAM_44_DMWIDTH/8-1:0] m_axis_bram_44_tstrb,
    output [C_OUTPUT_BRAM_44_DMWIDTH-1:0] m_axis_bram_44_tdata,
    input m_axis_bram_44_tready,
    input [C_OUTPUT_BRAM_44_ADDR_WIDTH-1:0] ap_bram_oarg_44_addr0,
    input [C_OUTPUT_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_din0,
    output [C_OUTPUT_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_dout0,
    input ap_bram_oarg_44_clk0,
    input ap_bram_oarg_44_rst0,
    input [C_OUTPUT_BRAM_44_WIDTH/8-1:0] ap_bram_oarg_44_we0,
    input ap_bram_oarg_44_en0,
    input [C_OUTPUT_BRAM_44_ADDR_WIDTH-1:0] ap_bram_oarg_44_addr1,
    input [C_OUTPUT_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_din1,
    output [C_OUTPUT_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_dout1,
    input ap_bram_oarg_44_clk1,
    input ap_bram_oarg_44_rst1,
    input [C_OUTPUT_BRAM_44_WIDTH/8-1:0] ap_bram_oarg_44_we1,
    input ap_bram_oarg_44_en1,
    //out AXI-Stream output interface 45
    output m_axis_bram_45_tlast,
    output m_axis_bram_45_tvalid,
    output [C_OUTPUT_BRAM_45_DMWIDTH/8-1:0] m_axis_bram_45_tkeep,
    output [C_OUTPUT_BRAM_45_DMWIDTH/8-1:0] m_axis_bram_45_tstrb,
    output [C_OUTPUT_BRAM_45_DMWIDTH-1:0] m_axis_bram_45_tdata,
    input m_axis_bram_45_tready,
    input [C_OUTPUT_BRAM_45_ADDR_WIDTH-1:0] ap_bram_oarg_45_addr0,
    input [C_OUTPUT_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_din0,
    output [C_OUTPUT_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_dout0,
    input ap_bram_oarg_45_clk0,
    input ap_bram_oarg_45_rst0,
    input [C_OUTPUT_BRAM_45_WIDTH/8-1:0] ap_bram_oarg_45_we0,
    input ap_bram_oarg_45_en0,
    input [C_OUTPUT_BRAM_45_ADDR_WIDTH-1:0] ap_bram_oarg_45_addr1,
    input [C_OUTPUT_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_din1,
    output [C_OUTPUT_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_dout1,
    input ap_bram_oarg_45_clk1,
    input ap_bram_oarg_45_rst1,
    input [C_OUTPUT_BRAM_45_WIDTH/8-1:0] ap_bram_oarg_45_we1,
    input ap_bram_oarg_45_en1,
    //out AXI-Stream output interface 46
    output m_axis_bram_46_tlast,
    output m_axis_bram_46_tvalid,
    output [C_OUTPUT_BRAM_46_DMWIDTH/8-1:0] m_axis_bram_46_tkeep,
    output [C_OUTPUT_BRAM_46_DMWIDTH/8-1:0] m_axis_bram_46_tstrb,
    output [C_OUTPUT_BRAM_46_DMWIDTH-1:0] m_axis_bram_46_tdata,
    input m_axis_bram_46_tready,
    input [C_OUTPUT_BRAM_46_ADDR_WIDTH-1:0] ap_bram_oarg_46_addr0,
    input [C_OUTPUT_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_din0,
    output [C_OUTPUT_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_dout0,
    input ap_bram_oarg_46_clk0,
    input ap_bram_oarg_46_rst0,
    input [C_OUTPUT_BRAM_46_WIDTH/8-1:0] ap_bram_oarg_46_we0,
    input ap_bram_oarg_46_en0,
    input [C_OUTPUT_BRAM_46_ADDR_WIDTH-1:0] ap_bram_oarg_46_addr1,
    input [C_OUTPUT_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_din1,
    output [C_OUTPUT_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_dout1,
    input ap_bram_oarg_46_clk1,
    input ap_bram_oarg_46_rst1,
    input [C_OUTPUT_BRAM_46_WIDTH/8-1:0] ap_bram_oarg_46_we1,
    input ap_bram_oarg_46_en1,
    //out AXI-Stream output interface 47
    output m_axis_bram_47_tlast,
    output m_axis_bram_47_tvalid,
    output [C_OUTPUT_BRAM_47_DMWIDTH/8-1:0] m_axis_bram_47_tkeep,
    output [C_OUTPUT_BRAM_47_DMWIDTH/8-1:0] m_axis_bram_47_tstrb,
    output [C_OUTPUT_BRAM_47_DMWIDTH-1:0] m_axis_bram_47_tdata,
    input m_axis_bram_47_tready,
    input [C_OUTPUT_BRAM_47_ADDR_WIDTH-1:0] ap_bram_oarg_47_addr0,
    input [C_OUTPUT_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_din0,
    output [C_OUTPUT_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_dout0,
    input ap_bram_oarg_47_clk0,
    input ap_bram_oarg_47_rst0,
    input [C_OUTPUT_BRAM_47_WIDTH/8-1:0] ap_bram_oarg_47_we0,
    input ap_bram_oarg_47_en0,
    input [C_OUTPUT_BRAM_47_ADDR_WIDTH-1:0] ap_bram_oarg_47_addr1,
    input [C_OUTPUT_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_din1,
    output [C_OUTPUT_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_dout1,
    input ap_bram_oarg_47_clk1,
    input ap_bram_oarg_47_rst1,
    input [C_OUTPUT_BRAM_47_WIDTH/8-1:0] ap_bram_oarg_47_we1,
    input ap_bram_oarg_47_en1,
    //out AXI-Stream output interface 48
    output m_axis_bram_48_tlast,
    output m_axis_bram_48_tvalid,
    output [C_OUTPUT_BRAM_48_DMWIDTH/8-1:0] m_axis_bram_48_tkeep,
    output [C_OUTPUT_BRAM_48_DMWIDTH/8-1:0] m_axis_bram_48_tstrb,
    output [C_OUTPUT_BRAM_48_DMWIDTH-1:0] m_axis_bram_48_tdata,
    input m_axis_bram_48_tready,
    input [C_OUTPUT_BRAM_48_ADDR_WIDTH-1:0] ap_bram_oarg_48_addr0,
    input [C_OUTPUT_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_din0,
    output [C_OUTPUT_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_dout0,
    input ap_bram_oarg_48_clk0,
    input ap_bram_oarg_48_rst0,
    input [C_OUTPUT_BRAM_48_WIDTH/8-1:0] ap_bram_oarg_48_we0,
    input ap_bram_oarg_48_en0,
    input [C_OUTPUT_BRAM_48_ADDR_WIDTH-1:0] ap_bram_oarg_48_addr1,
    input [C_OUTPUT_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_din1,
    output [C_OUTPUT_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_dout1,
    input ap_bram_oarg_48_clk1,
    input ap_bram_oarg_48_rst1,
    input [C_OUTPUT_BRAM_48_WIDTH/8-1:0] ap_bram_oarg_48_we1,
    input ap_bram_oarg_48_en1,
    //out AXI-Stream output interface 49
    output m_axis_bram_49_tlast,
    output m_axis_bram_49_tvalid,
    output [C_OUTPUT_BRAM_49_DMWIDTH/8-1:0] m_axis_bram_49_tkeep,
    output [C_OUTPUT_BRAM_49_DMWIDTH/8-1:0] m_axis_bram_49_tstrb,
    output [C_OUTPUT_BRAM_49_DMWIDTH-1:0] m_axis_bram_49_tdata,
    input m_axis_bram_49_tready,
    input [C_OUTPUT_BRAM_49_ADDR_WIDTH-1:0] ap_bram_oarg_49_addr0,
    input [C_OUTPUT_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_din0,
    output [C_OUTPUT_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_dout0,
    input ap_bram_oarg_49_clk0,
    input ap_bram_oarg_49_rst0,
    input [C_OUTPUT_BRAM_49_WIDTH/8-1:0] ap_bram_oarg_49_we0,
    input ap_bram_oarg_49_en0,
    input [C_OUTPUT_BRAM_49_ADDR_WIDTH-1:0] ap_bram_oarg_49_addr1,
    input [C_OUTPUT_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_din1,
    output [C_OUTPUT_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_dout1,
    input ap_bram_oarg_49_clk1,
    input ap_bram_oarg_49_rst1,
    input [C_OUTPUT_BRAM_49_WIDTH/8-1:0] ap_bram_oarg_49_we1,
    input ap_bram_oarg_49_en1,
    //out AXI-Stream output interface 50
    output m_axis_bram_50_tlast,
    output m_axis_bram_50_tvalid,
    output [C_OUTPUT_BRAM_50_DMWIDTH/8-1:0] m_axis_bram_50_tkeep,
    output [C_OUTPUT_BRAM_50_DMWIDTH/8-1:0] m_axis_bram_50_tstrb,
    output [C_OUTPUT_BRAM_50_DMWIDTH-1:0] m_axis_bram_50_tdata,
    input m_axis_bram_50_tready,
    input [C_OUTPUT_BRAM_50_ADDR_WIDTH-1:0] ap_bram_oarg_50_addr0,
    input [C_OUTPUT_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_din0,
    output [C_OUTPUT_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_dout0,
    input ap_bram_oarg_50_clk0,
    input ap_bram_oarg_50_rst0,
    input [C_OUTPUT_BRAM_50_WIDTH/8-1:0] ap_bram_oarg_50_we0,
    input ap_bram_oarg_50_en0,
    input [C_OUTPUT_BRAM_50_ADDR_WIDTH-1:0] ap_bram_oarg_50_addr1,
    input [C_OUTPUT_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_din1,
    output [C_OUTPUT_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_dout1,
    input ap_bram_oarg_50_clk1,
    input ap_bram_oarg_50_rst1,
    input [C_OUTPUT_BRAM_50_WIDTH/8-1:0] ap_bram_oarg_50_we1,
    input ap_bram_oarg_50_en1,
    //out AXI-Stream output interface 51
    output m_axis_bram_51_tlast,
    output m_axis_bram_51_tvalid,
    output [C_OUTPUT_BRAM_51_DMWIDTH/8-1:0] m_axis_bram_51_tkeep,
    output [C_OUTPUT_BRAM_51_DMWIDTH/8-1:0] m_axis_bram_51_tstrb,
    output [C_OUTPUT_BRAM_51_DMWIDTH-1:0] m_axis_bram_51_tdata,
    input m_axis_bram_51_tready,
    input [C_OUTPUT_BRAM_51_ADDR_WIDTH-1:0] ap_bram_oarg_51_addr0,
    input [C_OUTPUT_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_din0,
    output [C_OUTPUT_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_dout0,
    input ap_bram_oarg_51_clk0,
    input ap_bram_oarg_51_rst0,
    input [C_OUTPUT_BRAM_51_WIDTH/8-1:0] ap_bram_oarg_51_we0,
    input ap_bram_oarg_51_en0,
    input [C_OUTPUT_BRAM_51_ADDR_WIDTH-1:0] ap_bram_oarg_51_addr1,
    input [C_OUTPUT_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_din1,
    output [C_OUTPUT_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_dout1,
    input ap_bram_oarg_51_clk1,
    input ap_bram_oarg_51_rst1,
    input [C_OUTPUT_BRAM_51_WIDTH/8-1:0] ap_bram_oarg_51_we1,
    input ap_bram_oarg_51_en1,
    //out AXI-Stream output interface 52
    output m_axis_bram_52_tlast,
    output m_axis_bram_52_tvalid,
    output [C_OUTPUT_BRAM_52_DMWIDTH/8-1:0] m_axis_bram_52_tkeep,
    output [C_OUTPUT_BRAM_52_DMWIDTH/8-1:0] m_axis_bram_52_tstrb,
    output [C_OUTPUT_BRAM_52_DMWIDTH-1:0] m_axis_bram_52_tdata,
    input m_axis_bram_52_tready,
    input [C_OUTPUT_BRAM_52_ADDR_WIDTH-1:0] ap_bram_oarg_52_addr0,
    input [C_OUTPUT_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_din0,
    output [C_OUTPUT_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_dout0,
    input ap_bram_oarg_52_clk0,
    input ap_bram_oarg_52_rst0,
    input [C_OUTPUT_BRAM_52_WIDTH/8-1:0] ap_bram_oarg_52_we0,
    input ap_bram_oarg_52_en0,
    input [C_OUTPUT_BRAM_52_ADDR_WIDTH-1:0] ap_bram_oarg_52_addr1,
    input [C_OUTPUT_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_din1,
    output [C_OUTPUT_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_dout1,
    input ap_bram_oarg_52_clk1,
    input ap_bram_oarg_52_rst1,
    input [C_OUTPUT_BRAM_52_WIDTH/8-1:0] ap_bram_oarg_52_we1,
    input ap_bram_oarg_52_en1,
    //out AXI-Stream output interface 53
    output m_axis_bram_53_tlast,
    output m_axis_bram_53_tvalid,
    output [C_OUTPUT_BRAM_53_DMWIDTH/8-1:0] m_axis_bram_53_tkeep,
    output [C_OUTPUT_BRAM_53_DMWIDTH/8-1:0] m_axis_bram_53_tstrb,
    output [C_OUTPUT_BRAM_53_DMWIDTH-1:0] m_axis_bram_53_tdata,
    input m_axis_bram_53_tready,
    input [C_OUTPUT_BRAM_53_ADDR_WIDTH-1:0] ap_bram_oarg_53_addr0,
    input [C_OUTPUT_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_din0,
    output [C_OUTPUT_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_dout0,
    input ap_bram_oarg_53_clk0,
    input ap_bram_oarg_53_rst0,
    input [C_OUTPUT_BRAM_53_WIDTH/8-1:0] ap_bram_oarg_53_we0,
    input ap_bram_oarg_53_en0,
    input [C_OUTPUT_BRAM_53_ADDR_WIDTH-1:0] ap_bram_oarg_53_addr1,
    input [C_OUTPUT_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_din1,
    output [C_OUTPUT_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_dout1,
    input ap_bram_oarg_53_clk1,
    input ap_bram_oarg_53_rst1,
    input [C_OUTPUT_BRAM_53_WIDTH/8-1:0] ap_bram_oarg_53_we1,
    input ap_bram_oarg_53_en1,
    //out AXI-Stream output interface 54
    output m_axis_bram_54_tlast,
    output m_axis_bram_54_tvalid,
    output [C_OUTPUT_BRAM_54_DMWIDTH/8-1:0] m_axis_bram_54_tkeep,
    output [C_OUTPUT_BRAM_54_DMWIDTH/8-1:0] m_axis_bram_54_tstrb,
    output [C_OUTPUT_BRAM_54_DMWIDTH-1:0] m_axis_bram_54_tdata,
    input m_axis_bram_54_tready,
    input [C_OUTPUT_BRAM_54_ADDR_WIDTH-1:0] ap_bram_oarg_54_addr0,
    input [C_OUTPUT_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_din0,
    output [C_OUTPUT_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_dout0,
    input ap_bram_oarg_54_clk0,
    input ap_bram_oarg_54_rst0,
    input [C_OUTPUT_BRAM_54_WIDTH/8-1:0] ap_bram_oarg_54_we0,
    input ap_bram_oarg_54_en0,
    input [C_OUTPUT_BRAM_54_ADDR_WIDTH-1:0] ap_bram_oarg_54_addr1,
    input [C_OUTPUT_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_din1,
    output [C_OUTPUT_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_dout1,
    input ap_bram_oarg_54_clk1,
    input ap_bram_oarg_54_rst1,
    input [C_OUTPUT_BRAM_54_WIDTH/8-1:0] ap_bram_oarg_54_we1,
    input ap_bram_oarg_54_en1,
    //out AXI-Stream output interface 55
    output m_axis_bram_55_tlast,
    output m_axis_bram_55_tvalid,
    output [C_OUTPUT_BRAM_55_DMWIDTH/8-1:0] m_axis_bram_55_tkeep,
    output [C_OUTPUT_BRAM_55_DMWIDTH/8-1:0] m_axis_bram_55_tstrb,
    output [C_OUTPUT_BRAM_55_DMWIDTH-1:0] m_axis_bram_55_tdata,
    input m_axis_bram_55_tready,
    input [C_OUTPUT_BRAM_55_ADDR_WIDTH-1:0] ap_bram_oarg_55_addr0,
    input [C_OUTPUT_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_din0,
    output [C_OUTPUT_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_dout0,
    input ap_bram_oarg_55_clk0,
    input ap_bram_oarg_55_rst0,
    input [C_OUTPUT_BRAM_55_WIDTH/8-1:0] ap_bram_oarg_55_we0,
    input ap_bram_oarg_55_en0,
    input [C_OUTPUT_BRAM_55_ADDR_WIDTH-1:0] ap_bram_oarg_55_addr1,
    input [C_OUTPUT_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_din1,
    output [C_OUTPUT_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_dout1,
    input ap_bram_oarg_55_clk1,
    input ap_bram_oarg_55_rst1,
    input [C_OUTPUT_BRAM_55_WIDTH/8-1:0] ap_bram_oarg_55_we1,
    input ap_bram_oarg_55_en1,
    //out AXI-Stream output interface 56
    output m_axis_bram_56_tlast,
    output m_axis_bram_56_tvalid,
    output [C_OUTPUT_BRAM_56_DMWIDTH/8-1:0] m_axis_bram_56_tkeep,
    output [C_OUTPUT_BRAM_56_DMWIDTH/8-1:0] m_axis_bram_56_tstrb,
    output [C_OUTPUT_BRAM_56_DMWIDTH-1:0] m_axis_bram_56_tdata,
    input m_axis_bram_56_tready,
    input [C_OUTPUT_BRAM_56_ADDR_WIDTH-1:0] ap_bram_oarg_56_addr0,
    input [C_OUTPUT_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_din0,
    output [C_OUTPUT_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_dout0,
    input ap_bram_oarg_56_clk0,
    input ap_bram_oarg_56_rst0,
    input [C_OUTPUT_BRAM_56_WIDTH/8-1:0] ap_bram_oarg_56_we0,
    input ap_bram_oarg_56_en0,
    input [C_OUTPUT_BRAM_56_ADDR_WIDTH-1:0] ap_bram_oarg_56_addr1,
    input [C_OUTPUT_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_din1,
    output [C_OUTPUT_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_dout1,
    input ap_bram_oarg_56_clk1,
    input ap_bram_oarg_56_rst1,
    input [C_OUTPUT_BRAM_56_WIDTH/8-1:0] ap_bram_oarg_56_we1,
    input ap_bram_oarg_56_en1,
    //out AXI-Stream output interface 57
    output m_axis_bram_57_tlast,
    output m_axis_bram_57_tvalid,
    output [C_OUTPUT_BRAM_57_DMWIDTH/8-1:0] m_axis_bram_57_tkeep,
    output [C_OUTPUT_BRAM_57_DMWIDTH/8-1:0] m_axis_bram_57_tstrb,
    output [C_OUTPUT_BRAM_57_DMWIDTH-1:0] m_axis_bram_57_tdata,
    input m_axis_bram_57_tready,
    input [C_OUTPUT_BRAM_57_ADDR_WIDTH-1:0] ap_bram_oarg_57_addr0,
    input [C_OUTPUT_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_din0,
    output [C_OUTPUT_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_dout0,
    input ap_bram_oarg_57_clk0,
    input ap_bram_oarg_57_rst0,
    input [C_OUTPUT_BRAM_57_WIDTH/8-1:0] ap_bram_oarg_57_we0,
    input ap_bram_oarg_57_en0,
    input [C_OUTPUT_BRAM_57_ADDR_WIDTH-1:0] ap_bram_oarg_57_addr1,
    input [C_OUTPUT_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_din1,
    output [C_OUTPUT_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_dout1,
    input ap_bram_oarg_57_clk1,
    input ap_bram_oarg_57_rst1,
    input [C_OUTPUT_BRAM_57_WIDTH/8-1:0] ap_bram_oarg_57_we1,
    input ap_bram_oarg_57_en1,
    //out AXI-Stream output interface 58
    output m_axis_bram_58_tlast,
    output m_axis_bram_58_tvalid,
    output [C_OUTPUT_BRAM_58_DMWIDTH/8-1:0] m_axis_bram_58_tkeep,
    output [C_OUTPUT_BRAM_58_DMWIDTH/8-1:0] m_axis_bram_58_tstrb,
    output [C_OUTPUT_BRAM_58_DMWIDTH-1:0] m_axis_bram_58_tdata,
    input m_axis_bram_58_tready,
    input [C_OUTPUT_BRAM_58_ADDR_WIDTH-1:0] ap_bram_oarg_58_addr0,
    input [C_OUTPUT_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_din0,
    output [C_OUTPUT_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_dout0,
    input ap_bram_oarg_58_clk0,
    input ap_bram_oarg_58_rst0,
    input [C_OUTPUT_BRAM_58_WIDTH/8-1:0] ap_bram_oarg_58_we0,
    input ap_bram_oarg_58_en0,
    input [C_OUTPUT_BRAM_58_ADDR_WIDTH-1:0] ap_bram_oarg_58_addr1,
    input [C_OUTPUT_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_din1,
    output [C_OUTPUT_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_dout1,
    input ap_bram_oarg_58_clk1,
    input ap_bram_oarg_58_rst1,
    input [C_OUTPUT_BRAM_58_WIDTH/8-1:0] ap_bram_oarg_58_we1,
    input ap_bram_oarg_58_en1,
    //out AXI-Stream output interface 59
    output m_axis_bram_59_tlast,
    output m_axis_bram_59_tvalid,
    output [C_OUTPUT_BRAM_59_DMWIDTH/8-1:0] m_axis_bram_59_tkeep,
    output [C_OUTPUT_BRAM_59_DMWIDTH/8-1:0] m_axis_bram_59_tstrb,
    output [C_OUTPUT_BRAM_59_DMWIDTH-1:0] m_axis_bram_59_tdata,
    input m_axis_bram_59_tready,
    input [C_OUTPUT_BRAM_59_ADDR_WIDTH-1:0] ap_bram_oarg_59_addr0,
    input [C_OUTPUT_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_din0,
    output [C_OUTPUT_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_dout0,
    input ap_bram_oarg_59_clk0,
    input ap_bram_oarg_59_rst0,
    input [C_OUTPUT_BRAM_59_WIDTH/8-1:0] ap_bram_oarg_59_we0,
    input ap_bram_oarg_59_en0,
    input [C_OUTPUT_BRAM_59_ADDR_WIDTH-1:0] ap_bram_oarg_59_addr1,
    input [C_OUTPUT_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_din1,
    output [C_OUTPUT_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_dout1,
    input ap_bram_oarg_59_clk1,
    input ap_bram_oarg_59_rst1,
    input [C_OUTPUT_BRAM_59_WIDTH/8-1:0] ap_bram_oarg_59_we1,
    input ap_bram_oarg_59_en1,
    //out AXI-Stream output interface 60
    output m_axis_bram_60_tlast,
    output m_axis_bram_60_tvalid,
    output [C_OUTPUT_BRAM_60_DMWIDTH/8-1:0] m_axis_bram_60_tkeep,
    output [C_OUTPUT_BRAM_60_DMWIDTH/8-1:0] m_axis_bram_60_tstrb,
    output [C_OUTPUT_BRAM_60_DMWIDTH-1:0] m_axis_bram_60_tdata,
    input m_axis_bram_60_tready,
    input [C_OUTPUT_BRAM_60_ADDR_WIDTH-1:0] ap_bram_oarg_60_addr0,
    input [C_OUTPUT_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_din0,
    output [C_OUTPUT_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_dout0,
    input ap_bram_oarg_60_clk0,
    input ap_bram_oarg_60_rst0,
    input [C_OUTPUT_BRAM_60_WIDTH/8-1:0] ap_bram_oarg_60_we0,
    input ap_bram_oarg_60_en0,
    input [C_OUTPUT_BRAM_60_ADDR_WIDTH-1:0] ap_bram_oarg_60_addr1,
    input [C_OUTPUT_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_din1,
    output [C_OUTPUT_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_dout1,
    input ap_bram_oarg_60_clk1,
    input ap_bram_oarg_60_rst1,
    input [C_OUTPUT_BRAM_60_WIDTH/8-1:0] ap_bram_oarg_60_we1,
    input ap_bram_oarg_60_en1,
    //out AXI-Stream output interface 61
    output m_axis_bram_61_tlast,
    output m_axis_bram_61_tvalid,
    output [C_OUTPUT_BRAM_61_DMWIDTH/8-1:0] m_axis_bram_61_tkeep,
    output [C_OUTPUT_BRAM_61_DMWIDTH/8-1:0] m_axis_bram_61_tstrb,
    output [C_OUTPUT_BRAM_61_DMWIDTH-1:0] m_axis_bram_61_tdata,
    input m_axis_bram_61_tready,
    input [C_OUTPUT_BRAM_61_ADDR_WIDTH-1:0] ap_bram_oarg_61_addr0,
    input [C_OUTPUT_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_din0,
    output [C_OUTPUT_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_dout0,
    input ap_bram_oarg_61_clk0,
    input ap_bram_oarg_61_rst0,
    input [C_OUTPUT_BRAM_61_WIDTH/8-1:0] ap_bram_oarg_61_we0,
    input ap_bram_oarg_61_en0,
    input [C_OUTPUT_BRAM_61_ADDR_WIDTH-1:0] ap_bram_oarg_61_addr1,
    input [C_OUTPUT_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_din1,
    output [C_OUTPUT_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_dout1,
    input ap_bram_oarg_61_clk1,
    input ap_bram_oarg_61_rst1,
    input [C_OUTPUT_BRAM_61_WIDTH/8-1:0] ap_bram_oarg_61_we1,
    input ap_bram_oarg_61_en1,
    //out AXI-Stream output interface 62
    output m_axis_bram_62_tlast,
    output m_axis_bram_62_tvalid,
    output [C_OUTPUT_BRAM_62_DMWIDTH/8-1:0] m_axis_bram_62_tkeep,
    output [C_OUTPUT_BRAM_62_DMWIDTH/8-1:0] m_axis_bram_62_tstrb,
    output [C_OUTPUT_BRAM_62_DMWIDTH-1:0] m_axis_bram_62_tdata,
    input m_axis_bram_62_tready,
    input [C_OUTPUT_BRAM_62_ADDR_WIDTH-1:0] ap_bram_oarg_62_addr0,
    input [C_OUTPUT_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_din0,
    output [C_OUTPUT_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_dout0,
    input ap_bram_oarg_62_clk0,
    input ap_bram_oarg_62_rst0,
    input [C_OUTPUT_BRAM_62_WIDTH/8-1:0] ap_bram_oarg_62_we0,
    input ap_bram_oarg_62_en0,
    input [C_OUTPUT_BRAM_62_ADDR_WIDTH-1:0] ap_bram_oarg_62_addr1,
    input [C_OUTPUT_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_din1,
    output [C_OUTPUT_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_dout1,
    input ap_bram_oarg_62_clk1,
    input ap_bram_oarg_62_rst1,
    input [C_OUTPUT_BRAM_62_WIDTH/8-1:0] ap_bram_oarg_62_we1,
    input ap_bram_oarg_62_en1,
    //out AXI-Stream output interface 63
    output m_axis_bram_63_tlast,
    output m_axis_bram_63_tvalid,
    output [C_OUTPUT_BRAM_63_DMWIDTH/8-1:0] m_axis_bram_63_tkeep,
    output [C_OUTPUT_BRAM_63_DMWIDTH/8-1:0] m_axis_bram_63_tstrb,
    output [C_OUTPUT_BRAM_63_DMWIDTH-1:0] m_axis_bram_63_tdata,
    input m_axis_bram_63_tready,
    input [C_OUTPUT_BRAM_63_ADDR_WIDTH-1:0] ap_bram_oarg_63_addr0,
    input [C_OUTPUT_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_din0,
    output [C_OUTPUT_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_dout0,
    input ap_bram_oarg_63_clk0,
    input ap_bram_oarg_63_rst0,
    input [C_OUTPUT_BRAM_63_WIDTH/8-1:0] ap_bram_oarg_63_we0,
    input ap_bram_oarg_63_en0,
    input [C_OUTPUT_BRAM_63_ADDR_WIDTH-1:0] ap_bram_oarg_63_addr1,
    input [C_OUTPUT_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_din1,
    output [C_OUTPUT_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_dout1,
    input ap_bram_oarg_63_clk1,
    input ap_bram_oarg_63_rst1,
    input [C_OUTPUT_BRAM_63_WIDTH/8-1:0] ap_bram_oarg_63_we1,
    input ap_bram_oarg_63_en1,
    //out AXI-Stream output interface 64
    output m_axis_bram_64_tlast,
    output m_axis_bram_64_tvalid,
    output [C_OUTPUT_BRAM_64_DMWIDTH/8-1:0] m_axis_bram_64_tkeep,
    output [C_OUTPUT_BRAM_64_DMWIDTH/8-1:0] m_axis_bram_64_tstrb,
    output [C_OUTPUT_BRAM_64_DMWIDTH-1:0] m_axis_bram_64_tdata,
    input m_axis_bram_64_tready,
    input [C_OUTPUT_BRAM_64_ADDR_WIDTH-1:0] ap_bram_oarg_64_addr0,
    input [C_OUTPUT_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_din0,
    output [C_OUTPUT_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_dout0,
    input ap_bram_oarg_64_clk0,
    input ap_bram_oarg_64_rst0,
    input [C_OUTPUT_BRAM_64_WIDTH/8-1:0] ap_bram_oarg_64_we0,
    input ap_bram_oarg_64_en0,
    input [C_OUTPUT_BRAM_64_ADDR_WIDTH-1:0] ap_bram_oarg_64_addr1,
    input [C_OUTPUT_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_din1,
    output [C_OUTPUT_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_dout1,
    input ap_bram_oarg_64_clk1,
    input ap_bram_oarg_64_rst1,
    input [C_OUTPUT_BRAM_64_WIDTH/8-1:0] ap_bram_oarg_64_we1,
    input ap_bram_oarg_64_en1,
    //out AXI-Stream output interface 65
    output m_axis_bram_65_tlast,
    output m_axis_bram_65_tvalid,
    output [C_OUTPUT_BRAM_65_DMWIDTH/8-1:0] m_axis_bram_65_tkeep,
    output [C_OUTPUT_BRAM_65_DMWIDTH/8-1:0] m_axis_bram_65_tstrb,
    output [C_OUTPUT_BRAM_65_DMWIDTH-1:0] m_axis_bram_65_tdata,
    input m_axis_bram_65_tready,
    input [C_OUTPUT_BRAM_65_ADDR_WIDTH-1:0] ap_bram_oarg_65_addr0,
    input [C_OUTPUT_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_din0,
    output [C_OUTPUT_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_dout0,
    input ap_bram_oarg_65_clk0,
    input ap_bram_oarg_65_rst0,
    input [C_OUTPUT_BRAM_65_WIDTH/8-1:0] ap_bram_oarg_65_we0,
    input ap_bram_oarg_65_en0,
    input [C_OUTPUT_BRAM_65_ADDR_WIDTH-1:0] ap_bram_oarg_65_addr1,
    input [C_OUTPUT_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_din1,
    output [C_OUTPUT_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_dout1,
    input ap_bram_oarg_65_clk1,
    input ap_bram_oarg_65_rst1,
    input [C_OUTPUT_BRAM_65_WIDTH/8-1:0] ap_bram_oarg_65_we1,
    input ap_bram_oarg_65_en1,
    //out AXI-Stream output interface 66
    output m_axis_bram_66_tlast,
    output m_axis_bram_66_tvalid,
    output [C_OUTPUT_BRAM_66_DMWIDTH/8-1:0] m_axis_bram_66_tkeep,
    output [C_OUTPUT_BRAM_66_DMWIDTH/8-1:0] m_axis_bram_66_tstrb,
    output [C_OUTPUT_BRAM_66_DMWIDTH-1:0] m_axis_bram_66_tdata,
    input m_axis_bram_66_tready,
    input [C_OUTPUT_BRAM_66_ADDR_WIDTH-1:0] ap_bram_oarg_66_addr0,
    input [C_OUTPUT_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_din0,
    output [C_OUTPUT_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_dout0,
    input ap_bram_oarg_66_clk0,
    input ap_bram_oarg_66_rst0,
    input [C_OUTPUT_BRAM_66_WIDTH/8-1:0] ap_bram_oarg_66_we0,
    input ap_bram_oarg_66_en0,
    input [C_OUTPUT_BRAM_66_ADDR_WIDTH-1:0] ap_bram_oarg_66_addr1,
    input [C_OUTPUT_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_din1,
    output [C_OUTPUT_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_dout1,
    input ap_bram_oarg_66_clk1,
    input ap_bram_oarg_66_rst1,
    input [C_OUTPUT_BRAM_66_WIDTH/8-1:0] ap_bram_oarg_66_we1,
    input ap_bram_oarg_66_en1,
    //out AXI-Stream output interface 67
    output m_axis_bram_67_tlast,
    output m_axis_bram_67_tvalid,
    output [C_OUTPUT_BRAM_67_DMWIDTH/8-1:0] m_axis_bram_67_tkeep,
    output [C_OUTPUT_BRAM_67_DMWIDTH/8-1:0] m_axis_bram_67_tstrb,
    output [C_OUTPUT_BRAM_67_DMWIDTH-1:0] m_axis_bram_67_tdata,
    input m_axis_bram_67_tready,
    input [C_OUTPUT_BRAM_67_ADDR_WIDTH-1:0] ap_bram_oarg_67_addr0,
    input [C_OUTPUT_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_din0,
    output [C_OUTPUT_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_dout0,
    input ap_bram_oarg_67_clk0,
    input ap_bram_oarg_67_rst0,
    input [C_OUTPUT_BRAM_67_WIDTH/8-1:0] ap_bram_oarg_67_we0,
    input ap_bram_oarg_67_en0,
    input [C_OUTPUT_BRAM_67_ADDR_WIDTH-1:0] ap_bram_oarg_67_addr1,
    input [C_OUTPUT_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_din1,
    output [C_OUTPUT_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_dout1,
    input ap_bram_oarg_67_clk1,
    input ap_bram_oarg_67_rst1,
    input [C_OUTPUT_BRAM_67_WIDTH/8-1:0] ap_bram_oarg_67_we1,
    input ap_bram_oarg_67_en1,
    //out AXI-Stream output interface 68
    output m_axis_bram_68_tlast,
    output m_axis_bram_68_tvalid,
    output [C_OUTPUT_BRAM_68_DMWIDTH/8-1:0] m_axis_bram_68_tkeep,
    output [C_OUTPUT_BRAM_68_DMWIDTH/8-1:0] m_axis_bram_68_tstrb,
    output [C_OUTPUT_BRAM_68_DMWIDTH-1:0] m_axis_bram_68_tdata,
    input m_axis_bram_68_tready,
    input [C_OUTPUT_BRAM_68_ADDR_WIDTH-1:0] ap_bram_oarg_68_addr0,
    input [C_OUTPUT_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_din0,
    output [C_OUTPUT_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_dout0,
    input ap_bram_oarg_68_clk0,
    input ap_bram_oarg_68_rst0,
    input [C_OUTPUT_BRAM_68_WIDTH/8-1:0] ap_bram_oarg_68_we0,
    input ap_bram_oarg_68_en0,
    input [C_OUTPUT_BRAM_68_ADDR_WIDTH-1:0] ap_bram_oarg_68_addr1,
    input [C_OUTPUT_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_din1,
    output [C_OUTPUT_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_dout1,
    input ap_bram_oarg_68_clk1,
    input ap_bram_oarg_68_rst1,
    input [C_OUTPUT_BRAM_68_WIDTH/8-1:0] ap_bram_oarg_68_we1,
    input ap_bram_oarg_68_en1,
    //out AXI-Stream output interface 69
    output m_axis_bram_69_tlast,
    output m_axis_bram_69_tvalid,
    output [C_OUTPUT_BRAM_69_DMWIDTH/8-1:0] m_axis_bram_69_tkeep,
    output [C_OUTPUT_BRAM_69_DMWIDTH/8-1:0] m_axis_bram_69_tstrb,
    output [C_OUTPUT_BRAM_69_DMWIDTH-1:0] m_axis_bram_69_tdata,
    input m_axis_bram_69_tready,
    input [C_OUTPUT_BRAM_69_ADDR_WIDTH-1:0] ap_bram_oarg_69_addr0,
    input [C_OUTPUT_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_din0,
    output [C_OUTPUT_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_dout0,
    input ap_bram_oarg_69_clk0,
    input ap_bram_oarg_69_rst0,
    input [C_OUTPUT_BRAM_69_WIDTH/8-1:0] ap_bram_oarg_69_we0,
    input ap_bram_oarg_69_en0,
    input [C_OUTPUT_BRAM_69_ADDR_WIDTH-1:0] ap_bram_oarg_69_addr1,
    input [C_OUTPUT_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_din1,
    output [C_OUTPUT_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_dout1,
    input ap_bram_oarg_69_clk1,
    input ap_bram_oarg_69_rst1,
    input [C_OUTPUT_BRAM_69_WIDTH/8-1:0] ap_bram_oarg_69_we1,
    input ap_bram_oarg_69_en1,
    //out AXI-Stream output interface 70
    output m_axis_bram_70_tlast,
    output m_axis_bram_70_tvalid,
    output [C_OUTPUT_BRAM_70_DMWIDTH/8-1:0] m_axis_bram_70_tkeep,
    output [C_OUTPUT_BRAM_70_DMWIDTH/8-1:0] m_axis_bram_70_tstrb,
    output [C_OUTPUT_BRAM_70_DMWIDTH-1:0] m_axis_bram_70_tdata,
    input m_axis_bram_70_tready,
    input [C_OUTPUT_BRAM_70_ADDR_WIDTH-1:0] ap_bram_oarg_70_addr0,
    input [C_OUTPUT_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_din0,
    output [C_OUTPUT_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_dout0,
    input ap_bram_oarg_70_clk0,
    input ap_bram_oarg_70_rst0,
    input [C_OUTPUT_BRAM_70_WIDTH/8-1:0] ap_bram_oarg_70_we0,
    input ap_bram_oarg_70_en0,
    input [C_OUTPUT_BRAM_70_ADDR_WIDTH-1:0] ap_bram_oarg_70_addr1,
    input [C_OUTPUT_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_din1,
    output [C_OUTPUT_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_dout1,
    input ap_bram_oarg_70_clk1,
    input ap_bram_oarg_70_rst1,
    input [C_OUTPUT_BRAM_70_WIDTH/8-1:0] ap_bram_oarg_70_we1,
    input ap_bram_oarg_70_en1,
    //out AXI-Stream output interface 71
    output m_axis_bram_71_tlast,
    output m_axis_bram_71_tvalid,
    output [C_OUTPUT_BRAM_71_DMWIDTH/8-1:0] m_axis_bram_71_tkeep,
    output [C_OUTPUT_BRAM_71_DMWIDTH/8-1:0] m_axis_bram_71_tstrb,
    output [C_OUTPUT_BRAM_71_DMWIDTH-1:0] m_axis_bram_71_tdata,
    input m_axis_bram_71_tready,
    input [C_OUTPUT_BRAM_71_ADDR_WIDTH-1:0] ap_bram_oarg_71_addr0,
    input [C_OUTPUT_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_din0,
    output [C_OUTPUT_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_dout0,
    input ap_bram_oarg_71_clk0,
    input ap_bram_oarg_71_rst0,
    input [C_OUTPUT_BRAM_71_WIDTH/8-1:0] ap_bram_oarg_71_we0,
    input ap_bram_oarg_71_en0,
    input [C_OUTPUT_BRAM_71_ADDR_WIDTH-1:0] ap_bram_oarg_71_addr1,
    input [C_OUTPUT_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_din1,
    output [C_OUTPUT_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_dout1,
    input ap_bram_oarg_71_clk1,
    input ap_bram_oarg_71_rst1,
    input [C_OUTPUT_BRAM_71_WIDTH/8-1:0] ap_bram_oarg_71_we1,
    input ap_bram_oarg_71_en1,
    //out AXI-Stream output interface 72
    output m_axis_bram_72_tlast,
    output m_axis_bram_72_tvalid,
    output [C_OUTPUT_BRAM_72_DMWIDTH/8-1:0] m_axis_bram_72_tkeep,
    output [C_OUTPUT_BRAM_72_DMWIDTH/8-1:0] m_axis_bram_72_tstrb,
    output [C_OUTPUT_BRAM_72_DMWIDTH-1:0] m_axis_bram_72_tdata,
    input m_axis_bram_72_tready,
    input [C_OUTPUT_BRAM_72_ADDR_WIDTH-1:0] ap_bram_oarg_72_addr0,
    input [C_OUTPUT_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_din0,
    output [C_OUTPUT_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_dout0,
    input ap_bram_oarg_72_clk0,
    input ap_bram_oarg_72_rst0,
    input [C_OUTPUT_BRAM_72_WIDTH/8-1:0] ap_bram_oarg_72_we0,
    input ap_bram_oarg_72_en0,
    input [C_OUTPUT_BRAM_72_ADDR_WIDTH-1:0] ap_bram_oarg_72_addr1,
    input [C_OUTPUT_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_din1,
    output [C_OUTPUT_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_dout1,
    input ap_bram_oarg_72_clk1,
    input ap_bram_oarg_72_rst1,
    input [C_OUTPUT_BRAM_72_WIDTH/8-1:0] ap_bram_oarg_72_we1,
    input ap_bram_oarg_72_en1,
    //out AXI-Stream output interface 73
    output m_axis_bram_73_tlast,
    output m_axis_bram_73_tvalid,
    output [C_OUTPUT_BRAM_73_DMWIDTH/8-1:0] m_axis_bram_73_tkeep,
    output [C_OUTPUT_BRAM_73_DMWIDTH/8-1:0] m_axis_bram_73_tstrb,
    output [C_OUTPUT_BRAM_73_DMWIDTH-1:0] m_axis_bram_73_tdata,
    input m_axis_bram_73_tready,
    input [C_OUTPUT_BRAM_73_ADDR_WIDTH-1:0] ap_bram_oarg_73_addr0,
    input [C_OUTPUT_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_din0,
    output [C_OUTPUT_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_dout0,
    input ap_bram_oarg_73_clk0,
    input ap_bram_oarg_73_rst0,
    input [C_OUTPUT_BRAM_73_WIDTH/8-1:0] ap_bram_oarg_73_we0,
    input ap_bram_oarg_73_en0,
    input [C_OUTPUT_BRAM_73_ADDR_WIDTH-1:0] ap_bram_oarg_73_addr1,
    input [C_OUTPUT_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_din1,
    output [C_OUTPUT_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_dout1,
    input ap_bram_oarg_73_clk1,
    input ap_bram_oarg_73_rst1,
    input [C_OUTPUT_BRAM_73_WIDTH/8-1:0] ap_bram_oarg_73_we1,
    input ap_bram_oarg_73_en1,
    //out AXI-Stream output interface 74
    output m_axis_bram_74_tlast,
    output m_axis_bram_74_tvalid,
    output [C_OUTPUT_BRAM_74_DMWIDTH/8-1:0] m_axis_bram_74_tkeep,
    output [C_OUTPUT_BRAM_74_DMWIDTH/8-1:0] m_axis_bram_74_tstrb,
    output [C_OUTPUT_BRAM_74_DMWIDTH-1:0] m_axis_bram_74_tdata,
    input m_axis_bram_74_tready,
    input [C_OUTPUT_BRAM_74_ADDR_WIDTH-1:0] ap_bram_oarg_74_addr0,
    input [C_OUTPUT_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_din0,
    output [C_OUTPUT_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_dout0,
    input ap_bram_oarg_74_clk0,
    input ap_bram_oarg_74_rst0,
    input [C_OUTPUT_BRAM_74_WIDTH/8-1:0] ap_bram_oarg_74_we0,
    input ap_bram_oarg_74_en0,
    input [C_OUTPUT_BRAM_74_ADDR_WIDTH-1:0] ap_bram_oarg_74_addr1,
    input [C_OUTPUT_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_din1,
    output [C_OUTPUT_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_dout1,
    input ap_bram_oarg_74_clk1,
    input ap_bram_oarg_74_rst1,
    input [C_OUTPUT_BRAM_74_WIDTH/8-1:0] ap_bram_oarg_74_we1,
    input ap_bram_oarg_74_en1,
    //out AXI-Stream output interface 75
    output m_axis_bram_75_tlast,
    output m_axis_bram_75_tvalid,
    output [C_OUTPUT_BRAM_75_DMWIDTH/8-1:0] m_axis_bram_75_tkeep,
    output [C_OUTPUT_BRAM_75_DMWIDTH/8-1:0] m_axis_bram_75_tstrb,
    output [C_OUTPUT_BRAM_75_DMWIDTH-1:0] m_axis_bram_75_tdata,
    input m_axis_bram_75_tready,
    input [C_OUTPUT_BRAM_75_ADDR_WIDTH-1:0] ap_bram_oarg_75_addr0,
    input [C_OUTPUT_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_din0,
    output [C_OUTPUT_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_dout0,
    input ap_bram_oarg_75_clk0,
    input ap_bram_oarg_75_rst0,
    input [C_OUTPUT_BRAM_75_WIDTH/8-1:0] ap_bram_oarg_75_we0,
    input ap_bram_oarg_75_en0,
    input [C_OUTPUT_BRAM_75_ADDR_WIDTH-1:0] ap_bram_oarg_75_addr1,
    input [C_OUTPUT_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_din1,
    output [C_OUTPUT_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_dout1,
    input ap_bram_oarg_75_clk1,
    input ap_bram_oarg_75_rst1,
    input [C_OUTPUT_BRAM_75_WIDTH/8-1:0] ap_bram_oarg_75_we1,
    input ap_bram_oarg_75_en1,
    //out AXI-Stream output interface 76
    output m_axis_bram_76_tlast,
    output m_axis_bram_76_tvalid,
    output [C_OUTPUT_BRAM_76_DMWIDTH/8-1:0] m_axis_bram_76_tkeep,
    output [C_OUTPUT_BRAM_76_DMWIDTH/8-1:0] m_axis_bram_76_tstrb,
    output [C_OUTPUT_BRAM_76_DMWIDTH-1:0] m_axis_bram_76_tdata,
    input m_axis_bram_76_tready,
    input [C_OUTPUT_BRAM_76_ADDR_WIDTH-1:0] ap_bram_oarg_76_addr0,
    input [C_OUTPUT_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_din0,
    output [C_OUTPUT_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_dout0,
    input ap_bram_oarg_76_clk0,
    input ap_bram_oarg_76_rst0,
    input [C_OUTPUT_BRAM_76_WIDTH/8-1:0] ap_bram_oarg_76_we0,
    input ap_bram_oarg_76_en0,
    input [C_OUTPUT_BRAM_76_ADDR_WIDTH-1:0] ap_bram_oarg_76_addr1,
    input [C_OUTPUT_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_din1,
    output [C_OUTPUT_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_dout1,
    input ap_bram_oarg_76_clk1,
    input ap_bram_oarg_76_rst1,
    input [C_OUTPUT_BRAM_76_WIDTH/8-1:0] ap_bram_oarg_76_we1,
    input ap_bram_oarg_76_en1,
    //out AXI-Stream output interface 77
    output m_axis_bram_77_tlast,
    output m_axis_bram_77_tvalid,
    output [C_OUTPUT_BRAM_77_DMWIDTH/8-1:0] m_axis_bram_77_tkeep,
    output [C_OUTPUT_BRAM_77_DMWIDTH/8-1:0] m_axis_bram_77_tstrb,
    output [C_OUTPUT_BRAM_77_DMWIDTH-1:0] m_axis_bram_77_tdata,
    input m_axis_bram_77_tready,
    input [C_OUTPUT_BRAM_77_ADDR_WIDTH-1:0] ap_bram_oarg_77_addr0,
    input [C_OUTPUT_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_din0,
    output [C_OUTPUT_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_dout0,
    input ap_bram_oarg_77_clk0,
    input ap_bram_oarg_77_rst0,
    input [C_OUTPUT_BRAM_77_WIDTH/8-1:0] ap_bram_oarg_77_we0,
    input ap_bram_oarg_77_en0,
    input [C_OUTPUT_BRAM_77_ADDR_WIDTH-1:0] ap_bram_oarg_77_addr1,
    input [C_OUTPUT_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_din1,
    output [C_OUTPUT_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_dout1,
    input ap_bram_oarg_77_clk1,
    input ap_bram_oarg_77_rst1,
    input [C_OUTPUT_BRAM_77_WIDTH/8-1:0] ap_bram_oarg_77_we1,
    input ap_bram_oarg_77_en1,
    //out AXI-Stream output interface 78
    output m_axis_bram_78_tlast,
    output m_axis_bram_78_tvalid,
    output [C_OUTPUT_BRAM_78_DMWIDTH/8-1:0] m_axis_bram_78_tkeep,
    output [C_OUTPUT_BRAM_78_DMWIDTH/8-1:0] m_axis_bram_78_tstrb,
    output [C_OUTPUT_BRAM_78_DMWIDTH-1:0] m_axis_bram_78_tdata,
    input m_axis_bram_78_tready,
    input [C_OUTPUT_BRAM_78_ADDR_WIDTH-1:0] ap_bram_oarg_78_addr0,
    input [C_OUTPUT_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_din0,
    output [C_OUTPUT_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_dout0,
    input ap_bram_oarg_78_clk0,
    input ap_bram_oarg_78_rst0,
    input [C_OUTPUT_BRAM_78_WIDTH/8-1:0] ap_bram_oarg_78_we0,
    input ap_bram_oarg_78_en0,
    input [C_OUTPUT_BRAM_78_ADDR_WIDTH-1:0] ap_bram_oarg_78_addr1,
    input [C_OUTPUT_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_din1,
    output [C_OUTPUT_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_dout1,
    input ap_bram_oarg_78_clk1,
    input ap_bram_oarg_78_rst1,
    input [C_OUTPUT_BRAM_78_WIDTH/8-1:0] ap_bram_oarg_78_we1,
    input ap_bram_oarg_78_en1,
    //out AXI-Stream output interface 79
    output m_axis_bram_79_tlast,
    output m_axis_bram_79_tvalid,
    output [C_OUTPUT_BRAM_79_DMWIDTH/8-1:0] m_axis_bram_79_tkeep,
    output [C_OUTPUT_BRAM_79_DMWIDTH/8-1:0] m_axis_bram_79_tstrb,
    output [C_OUTPUT_BRAM_79_DMWIDTH-1:0] m_axis_bram_79_tdata,
    input m_axis_bram_79_tready,
    input [C_OUTPUT_BRAM_79_ADDR_WIDTH-1:0] ap_bram_oarg_79_addr0,
    input [C_OUTPUT_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_din0,
    output [C_OUTPUT_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_dout0,
    input ap_bram_oarg_79_clk0,
    input ap_bram_oarg_79_rst0,
    input [C_OUTPUT_BRAM_79_WIDTH/8-1:0] ap_bram_oarg_79_we0,
    input ap_bram_oarg_79_en0,
    input [C_OUTPUT_BRAM_79_ADDR_WIDTH-1:0] ap_bram_oarg_79_addr1,
    input [C_OUTPUT_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_din1,
    output [C_OUTPUT_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_dout1,
    input ap_bram_oarg_79_clk1,
    input ap_bram_oarg_79_rst1,
    input [C_OUTPUT_BRAM_79_WIDTH/8-1:0] ap_bram_oarg_79_we1,
    input ap_bram_oarg_79_en1,
    //out AXI-Stream output interface 80
    output m_axis_bram_80_tlast,
    output m_axis_bram_80_tvalid,
    output [C_OUTPUT_BRAM_80_DMWIDTH/8-1:0] m_axis_bram_80_tkeep,
    output [C_OUTPUT_BRAM_80_DMWIDTH/8-1:0] m_axis_bram_80_tstrb,
    output [C_OUTPUT_BRAM_80_DMWIDTH-1:0] m_axis_bram_80_tdata,
    input m_axis_bram_80_tready,
    input [C_OUTPUT_BRAM_80_ADDR_WIDTH-1:0] ap_bram_oarg_80_addr0,
    input [C_OUTPUT_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_din0,
    output [C_OUTPUT_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_dout0,
    input ap_bram_oarg_80_clk0,
    input ap_bram_oarg_80_rst0,
    input [C_OUTPUT_BRAM_80_WIDTH/8-1:0] ap_bram_oarg_80_we0,
    input ap_bram_oarg_80_en0,
    input [C_OUTPUT_BRAM_80_ADDR_WIDTH-1:0] ap_bram_oarg_80_addr1,
    input [C_OUTPUT_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_din1,
    output [C_OUTPUT_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_dout1,
    input ap_bram_oarg_80_clk1,
    input ap_bram_oarg_80_rst1,
    input [C_OUTPUT_BRAM_80_WIDTH/8-1:0] ap_bram_oarg_80_we1,
    input ap_bram_oarg_80_en1,
    //out AXI-Stream output interface 81
    output m_axis_bram_81_tlast,
    output m_axis_bram_81_tvalid,
    output [C_OUTPUT_BRAM_81_DMWIDTH/8-1:0] m_axis_bram_81_tkeep,
    output [C_OUTPUT_BRAM_81_DMWIDTH/8-1:0] m_axis_bram_81_tstrb,
    output [C_OUTPUT_BRAM_81_DMWIDTH-1:0] m_axis_bram_81_tdata,
    input m_axis_bram_81_tready,
    input [C_OUTPUT_BRAM_81_ADDR_WIDTH-1:0] ap_bram_oarg_81_addr0,
    input [C_OUTPUT_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_din0,
    output [C_OUTPUT_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_dout0,
    input ap_bram_oarg_81_clk0,
    input ap_bram_oarg_81_rst0,
    input [C_OUTPUT_BRAM_81_WIDTH/8-1:0] ap_bram_oarg_81_we0,
    input ap_bram_oarg_81_en0,
    input [C_OUTPUT_BRAM_81_ADDR_WIDTH-1:0] ap_bram_oarg_81_addr1,
    input [C_OUTPUT_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_din1,
    output [C_OUTPUT_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_dout1,
    input ap_bram_oarg_81_clk1,
    input ap_bram_oarg_81_rst1,
    input [C_OUTPUT_BRAM_81_WIDTH/8-1:0] ap_bram_oarg_81_we1,
    input ap_bram_oarg_81_en1,
    //out AXI-Stream output interface 82
    output m_axis_bram_82_tlast,
    output m_axis_bram_82_tvalid,
    output [C_OUTPUT_BRAM_82_DMWIDTH/8-1:0] m_axis_bram_82_tkeep,
    output [C_OUTPUT_BRAM_82_DMWIDTH/8-1:0] m_axis_bram_82_tstrb,
    output [C_OUTPUT_BRAM_82_DMWIDTH-1:0] m_axis_bram_82_tdata,
    input m_axis_bram_82_tready,
    input [C_OUTPUT_BRAM_82_ADDR_WIDTH-1:0] ap_bram_oarg_82_addr0,
    input [C_OUTPUT_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_din0,
    output [C_OUTPUT_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_dout0,
    input ap_bram_oarg_82_clk0,
    input ap_bram_oarg_82_rst0,
    input [C_OUTPUT_BRAM_82_WIDTH/8-1:0] ap_bram_oarg_82_we0,
    input ap_bram_oarg_82_en0,
    input [C_OUTPUT_BRAM_82_ADDR_WIDTH-1:0] ap_bram_oarg_82_addr1,
    input [C_OUTPUT_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_din1,
    output [C_OUTPUT_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_dout1,
    input ap_bram_oarg_82_clk1,
    input ap_bram_oarg_82_rst1,
    input [C_OUTPUT_BRAM_82_WIDTH/8-1:0] ap_bram_oarg_82_we1,
    input ap_bram_oarg_82_en1,
    //out AXI-Stream output interface 83
    output m_axis_bram_83_tlast,
    output m_axis_bram_83_tvalid,
    output [C_OUTPUT_BRAM_83_DMWIDTH/8-1:0] m_axis_bram_83_tkeep,
    output [C_OUTPUT_BRAM_83_DMWIDTH/8-1:0] m_axis_bram_83_tstrb,
    output [C_OUTPUT_BRAM_83_DMWIDTH-1:0] m_axis_bram_83_tdata,
    input m_axis_bram_83_tready,
    input [C_OUTPUT_BRAM_83_ADDR_WIDTH-1:0] ap_bram_oarg_83_addr0,
    input [C_OUTPUT_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_din0,
    output [C_OUTPUT_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_dout0,
    input ap_bram_oarg_83_clk0,
    input ap_bram_oarg_83_rst0,
    input [C_OUTPUT_BRAM_83_WIDTH/8-1:0] ap_bram_oarg_83_we0,
    input ap_bram_oarg_83_en0,
    input [C_OUTPUT_BRAM_83_ADDR_WIDTH-1:0] ap_bram_oarg_83_addr1,
    input [C_OUTPUT_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_din1,
    output [C_OUTPUT_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_dout1,
    input ap_bram_oarg_83_clk1,
    input ap_bram_oarg_83_rst1,
    input [C_OUTPUT_BRAM_83_WIDTH/8-1:0] ap_bram_oarg_83_we1,
    input ap_bram_oarg_83_en1,
    //out AXI-Stream output interface 84
    output m_axis_bram_84_tlast,
    output m_axis_bram_84_tvalid,
    output [C_OUTPUT_BRAM_84_DMWIDTH/8-1:0] m_axis_bram_84_tkeep,
    output [C_OUTPUT_BRAM_84_DMWIDTH/8-1:0] m_axis_bram_84_tstrb,
    output [C_OUTPUT_BRAM_84_DMWIDTH-1:0] m_axis_bram_84_tdata,
    input m_axis_bram_84_tready,
    input [C_OUTPUT_BRAM_84_ADDR_WIDTH-1:0] ap_bram_oarg_84_addr0,
    input [C_OUTPUT_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_din0,
    output [C_OUTPUT_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_dout0,
    input ap_bram_oarg_84_clk0,
    input ap_bram_oarg_84_rst0,
    input [C_OUTPUT_BRAM_84_WIDTH/8-1:0] ap_bram_oarg_84_we0,
    input ap_bram_oarg_84_en0,
    input [C_OUTPUT_BRAM_84_ADDR_WIDTH-1:0] ap_bram_oarg_84_addr1,
    input [C_OUTPUT_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_din1,
    output [C_OUTPUT_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_dout1,
    input ap_bram_oarg_84_clk1,
    input ap_bram_oarg_84_rst1,
    input [C_OUTPUT_BRAM_84_WIDTH/8-1:0] ap_bram_oarg_84_we1,
    input ap_bram_oarg_84_en1,
    //out AXI-Stream output interface 85
    output m_axis_bram_85_tlast,
    output m_axis_bram_85_tvalid,
    output [C_OUTPUT_BRAM_85_DMWIDTH/8-1:0] m_axis_bram_85_tkeep,
    output [C_OUTPUT_BRAM_85_DMWIDTH/8-1:0] m_axis_bram_85_tstrb,
    output [C_OUTPUT_BRAM_85_DMWIDTH-1:0] m_axis_bram_85_tdata,
    input m_axis_bram_85_tready,
    input [C_OUTPUT_BRAM_85_ADDR_WIDTH-1:0] ap_bram_oarg_85_addr0,
    input [C_OUTPUT_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_din0,
    output [C_OUTPUT_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_dout0,
    input ap_bram_oarg_85_clk0,
    input ap_bram_oarg_85_rst0,
    input [C_OUTPUT_BRAM_85_WIDTH/8-1:0] ap_bram_oarg_85_we0,
    input ap_bram_oarg_85_en0,
    input [C_OUTPUT_BRAM_85_ADDR_WIDTH-1:0] ap_bram_oarg_85_addr1,
    input [C_OUTPUT_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_din1,
    output [C_OUTPUT_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_dout1,
    input ap_bram_oarg_85_clk1,
    input ap_bram_oarg_85_rst1,
    input [C_OUTPUT_BRAM_85_WIDTH/8-1:0] ap_bram_oarg_85_we1,
    input ap_bram_oarg_85_en1,
    //out AXI-Stream output interface 86
    output m_axis_bram_86_tlast,
    output m_axis_bram_86_tvalid,
    output [C_OUTPUT_BRAM_86_DMWIDTH/8-1:0] m_axis_bram_86_tkeep,
    output [C_OUTPUT_BRAM_86_DMWIDTH/8-1:0] m_axis_bram_86_tstrb,
    output [C_OUTPUT_BRAM_86_DMWIDTH-1:0] m_axis_bram_86_tdata,
    input m_axis_bram_86_tready,
    input [C_OUTPUT_BRAM_86_ADDR_WIDTH-1:0] ap_bram_oarg_86_addr0,
    input [C_OUTPUT_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_din0,
    output [C_OUTPUT_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_dout0,
    input ap_bram_oarg_86_clk0,
    input ap_bram_oarg_86_rst0,
    input [C_OUTPUT_BRAM_86_WIDTH/8-1:0] ap_bram_oarg_86_we0,
    input ap_bram_oarg_86_en0,
    input [C_OUTPUT_BRAM_86_ADDR_WIDTH-1:0] ap_bram_oarg_86_addr1,
    input [C_OUTPUT_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_din1,
    output [C_OUTPUT_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_dout1,
    input ap_bram_oarg_86_clk1,
    input ap_bram_oarg_86_rst1,
    input [C_OUTPUT_BRAM_86_WIDTH/8-1:0] ap_bram_oarg_86_we1,
    input ap_bram_oarg_86_en1,
    //out AXI-Stream output interface 87
    output m_axis_bram_87_tlast,
    output m_axis_bram_87_tvalid,
    output [C_OUTPUT_BRAM_87_DMWIDTH/8-1:0] m_axis_bram_87_tkeep,
    output [C_OUTPUT_BRAM_87_DMWIDTH/8-1:0] m_axis_bram_87_tstrb,
    output [C_OUTPUT_BRAM_87_DMWIDTH-1:0] m_axis_bram_87_tdata,
    input m_axis_bram_87_tready,
    input [C_OUTPUT_BRAM_87_ADDR_WIDTH-1:0] ap_bram_oarg_87_addr0,
    input [C_OUTPUT_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_din0,
    output [C_OUTPUT_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_dout0,
    input ap_bram_oarg_87_clk0,
    input ap_bram_oarg_87_rst0,
    input [C_OUTPUT_BRAM_87_WIDTH/8-1:0] ap_bram_oarg_87_we0,
    input ap_bram_oarg_87_en0,
    input [C_OUTPUT_BRAM_87_ADDR_WIDTH-1:0] ap_bram_oarg_87_addr1,
    input [C_OUTPUT_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_din1,
    output [C_OUTPUT_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_dout1,
    input ap_bram_oarg_87_clk1,
    input ap_bram_oarg_87_rst1,
    input [C_OUTPUT_BRAM_87_WIDTH/8-1:0] ap_bram_oarg_87_we1,
    input ap_bram_oarg_87_en1,
    //out AXI-Stream output interface 88
    output m_axis_bram_88_tlast,
    output m_axis_bram_88_tvalid,
    output [C_OUTPUT_BRAM_88_DMWIDTH/8-1:0] m_axis_bram_88_tkeep,
    output [C_OUTPUT_BRAM_88_DMWIDTH/8-1:0] m_axis_bram_88_tstrb,
    output [C_OUTPUT_BRAM_88_DMWIDTH-1:0] m_axis_bram_88_tdata,
    input m_axis_bram_88_tready,
    input [C_OUTPUT_BRAM_88_ADDR_WIDTH-1:0] ap_bram_oarg_88_addr0,
    input [C_OUTPUT_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_din0,
    output [C_OUTPUT_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_dout0,
    input ap_bram_oarg_88_clk0,
    input ap_bram_oarg_88_rst0,
    input [C_OUTPUT_BRAM_88_WIDTH/8-1:0] ap_bram_oarg_88_we0,
    input ap_bram_oarg_88_en0,
    input [C_OUTPUT_BRAM_88_ADDR_WIDTH-1:0] ap_bram_oarg_88_addr1,
    input [C_OUTPUT_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_din1,
    output [C_OUTPUT_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_dout1,
    input ap_bram_oarg_88_clk1,
    input ap_bram_oarg_88_rst1,
    input [C_OUTPUT_BRAM_88_WIDTH/8-1:0] ap_bram_oarg_88_we1,
    input ap_bram_oarg_88_en1,
    //out AXI-Stream output interface 89
    output m_axis_bram_89_tlast,
    output m_axis_bram_89_tvalid,
    output [C_OUTPUT_BRAM_89_DMWIDTH/8-1:0] m_axis_bram_89_tkeep,
    output [C_OUTPUT_BRAM_89_DMWIDTH/8-1:0] m_axis_bram_89_tstrb,
    output [C_OUTPUT_BRAM_89_DMWIDTH-1:0] m_axis_bram_89_tdata,
    input m_axis_bram_89_tready,
    input [C_OUTPUT_BRAM_89_ADDR_WIDTH-1:0] ap_bram_oarg_89_addr0,
    input [C_OUTPUT_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_din0,
    output [C_OUTPUT_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_dout0,
    input ap_bram_oarg_89_clk0,
    input ap_bram_oarg_89_rst0,
    input [C_OUTPUT_BRAM_89_WIDTH/8-1:0] ap_bram_oarg_89_we0,
    input ap_bram_oarg_89_en0,
    input [C_OUTPUT_BRAM_89_ADDR_WIDTH-1:0] ap_bram_oarg_89_addr1,
    input [C_OUTPUT_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_din1,
    output [C_OUTPUT_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_dout1,
    input ap_bram_oarg_89_clk1,
    input ap_bram_oarg_89_rst1,
    input [C_OUTPUT_BRAM_89_WIDTH/8-1:0] ap_bram_oarg_89_we1,
    input ap_bram_oarg_89_en1,
    //out AXI-Stream output interface 90
    output m_axis_bram_90_tlast,
    output m_axis_bram_90_tvalid,
    output [C_OUTPUT_BRAM_90_DMWIDTH/8-1:0] m_axis_bram_90_tkeep,
    output [C_OUTPUT_BRAM_90_DMWIDTH/8-1:0] m_axis_bram_90_tstrb,
    output [C_OUTPUT_BRAM_90_DMWIDTH-1:0] m_axis_bram_90_tdata,
    input m_axis_bram_90_tready,
    input [C_OUTPUT_BRAM_90_ADDR_WIDTH-1:0] ap_bram_oarg_90_addr0,
    input [C_OUTPUT_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_din0,
    output [C_OUTPUT_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_dout0,
    input ap_bram_oarg_90_clk0,
    input ap_bram_oarg_90_rst0,
    input [C_OUTPUT_BRAM_90_WIDTH/8-1:0] ap_bram_oarg_90_we0,
    input ap_bram_oarg_90_en0,
    input [C_OUTPUT_BRAM_90_ADDR_WIDTH-1:0] ap_bram_oarg_90_addr1,
    input [C_OUTPUT_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_din1,
    output [C_OUTPUT_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_dout1,
    input ap_bram_oarg_90_clk1,
    input ap_bram_oarg_90_rst1,
    input [C_OUTPUT_BRAM_90_WIDTH/8-1:0] ap_bram_oarg_90_we1,
    input ap_bram_oarg_90_en1,
    //out AXI-Stream output interface 91
    output m_axis_bram_91_tlast,
    output m_axis_bram_91_tvalid,
    output [C_OUTPUT_BRAM_91_DMWIDTH/8-1:0] m_axis_bram_91_tkeep,
    output [C_OUTPUT_BRAM_91_DMWIDTH/8-1:0] m_axis_bram_91_tstrb,
    output [C_OUTPUT_BRAM_91_DMWIDTH-1:0] m_axis_bram_91_tdata,
    input m_axis_bram_91_tready,
    input [C_OUTPUT_BRAM_91_ADDR_WIDTH-1:0] ap_bram_oarg_91_addr0,
    input [C_OUTPUT_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_din0,
    output [C_OUTPUT_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_dout0,
    input ap_bram_oarg_91_clk0,
    input ap_bram_oarg_91_rst0,
    input [C_OUTPUT_BRAM_91_WIDTH/8-1:0] ap_bram_oarg_91_we0,
    input ap_bram_oarg_91_en0,
    input [C_OUTPUT_BRAM_91_ADDR_WIDTH-1:0] ap_bram_oarg_91_addr1,
    input [C_OUTPUT_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_din1,
    output [C_OUTPUT_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_dout1,
    input ap_bram_oarg_91_clk1,
    input ap_bram_oarg_91_rst1,
    input [C_OUTPUT_BRAM_91_WIDTH/8-1:0] ap_bram_oarg_91_we1,
    input ap_bram_oarg_91_en1,
    //out AXI-Stream output interface 92
    output m_axis_bram_92_tlast,
    output m_axis_bram_92_tvalid,
    output [C_OUTPUT_BRAM_92_DMWIDTH/8-1:0] m_axis_bram_92_tkeep,
    output [C_OUTPUT_BRAM_92_DMWIDTH/8-1:0] m_axis_bram_92_tstrb,
    output [C_OUTPUT_BRAM_92_DMWIDTH-1:0] m_axis_bram_92_tdata,
    input m_axis_bram_92_tready,
    input [C_OUTPUT_BRAM_92_ADDR_WIDTH-1:0] ap_bram_oarg_92_addr0,
    input [C_OUTPUT_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_din0,
    output [C_OUTPUT_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_dout0,
    input ap_bram_oarg_92_clk0,
    input ap_bram_oarg_92_rst0,
    input [C_OUTPUT_BRAM_92_WIDTH/8-1:0] ap_bram_oarg_92_we0,
    input ap_bram_oarg_92_en0,
    input [C_OUTPUT_BRAM_92_ADDR_WIDTH-1:0] ap_bram_oarg_92_addr1,
    input [C_OUTPUT_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_din1,
    output [C_OUTPUT_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_dout1,
    input ap_bram_oarg_92_clk1,
    input ap_bram_oarg_92_rst1,
    input [C_OUTPUT_BRAM_92_WIDTH/8-1:0] ap_bram_oarg_92_we1,
    input ap_bram_oarg_92_en1,
    //out AXI-Stream output interface 93
    output m_axis_bram_93_tlast,
    output m_axis_bram_93_tvalid,
    output [C_OUTPUT_BRAM_93_DMWIDTH/8-1:0] m_axis_bram_93_tkeep,
    output [C_OUTPUT_BRAM_93_DMWIDTH/8-1:0] m_axis_bram_93_tstrb,
    output [C_OUTPUT_BRAM_93_DMWIDTH-1:0] m_axis_bram_93_tdata,
    input m_axis_bram_93_tready,
    input [C_OUTPUT_BRAM_93_ADDR_WIDTH-1:0] ap_bram_oarg_93_addr0,
    input [C_OUTPUT_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_din0,
    output [C_OUTPUT_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_dout0,
    input ap_bram_oarg_93_clk0,
    input ap_bram_oarg_93_rst0,
    input [C_OUTPUT_BRAM_93_WIDTH/8-1:0] ap_bram_oarg_93_we0,
    input ap_bram_oarg_93_en0,
    input [C_OUTPUT_BRAM_93_ADDR_WIDTH-1:0] ap_bram_oarg_93_addr1,
    input [C_OUTPUT_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_din1,
    output [C_OUTPUT_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_dout1,
    input ap_bram_oarg_93_clk1,
    input ap_bram_oarg_93_rst1,
    input [C_OUTPUT_BRAM_93_WIDTH/8-1:0] ap_bram_oarg_93_we1,
    input ap_bram_oarg_93_en1,
    //out AXI-Stream output interface 94
    output m_axis_bram_94_tlast,
    output m_axis_bram_94_tvalid,
    output [C_OUTPUT_BRAM_94_DMWIDTH/8-1:0] m_axis_bram_94_tkeep,
    output [C_OUTPUT_BRAM_94_DMWIDTH/8-1:0] m_axis_bram_94_tstrb,
    output [C_OUTPUT_BRAM_94_DMWIDTH-1:0] m_axis_bram_94_tdata,
    input m_axis_bram_94_tready,
    input [C_OUTPUT_BRAM_94_ADDR_WIDTH-1:0] ap_bram_oarg_94_addr0,
    input [C_OUTPUT_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_din0,
    output [C_OUTPUT_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_dout0,
    input ap_bram_oarg_94_clk0,
    input ap_bram_oarg_94_rst0,
    input [C_OUTPUT_BRAM_94_WIDTH/8-1:0] ap_bram_oarg_94_we0,
    input ap_bram_oarg_94_en0,
    input [C_OUTPUT_BRAM_94_ADDR_WIDTH-1:0] ap_bram_oarg_94_addr1,
    input [C_OUTPUT_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_din1,
    output [C_OUTPUT_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_dout1,
    input ap_bram_oarg_94_clk1,
    input ap_bram_oarg_94_rst1,
    input [C_OUTPUT_BRAM_94_WIDTH/8-1:0] ap_bram_oarg_94_we1,
    input ap_bram_oarg_94_en1,
    //out AXI-Stream output interface 95
    output m_axis_bram_95_tlast,
    output m_axis_bram_95_tvalid,
    output [C_OUTPUT_BRAM_95_DMWIDTH/8-1:0] m_axis_bram_95_tkeep,
    output [C_OUTPUT_BRAM_95_DMWIDTH/8-1:0] m_axis_bram_95_tstrb,
    output [C_OUTPUT_BRAM_95_DMWIDTH-1:0] m_axis_bram_95_tdata,
    input m_axis_bram_95_tready,
    input [C_OUTPUT_BRAM_95_ADDR_WIDTH-1:0] ap_bram_oarg_95_addr0,
    input [C_OUTPUT_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_din0,
    output [C_OUTPUT_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_dout0,
    input ap_bram_oarg_95_clk0,
    input ap_bram_oarg_95_rst0,
    input [C_OUTPUT_BRAM_95_WIDTH/8-1:0] ap_bram_oarg_95_we0,
    input ap_bram_oarg_95_en0,
    input [C_OUTPUT_BRAM_95_ADDR_WIDTH-1:0] ap_bram_oarg_95_addr1,
    input [C_OUTPUT_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_din1,
    output [C_OUTPUT_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_dout1,
    input ap_bram_oarg_95_clk1,
    input ap_bram_oarg_95_rst1,
    input [C_OUTPUT_BRAM_95_WIDTH/8-1:0] ap_bram_oarg_95_we1,
    input ap_bram_oarg_95_en1,
    //out AXI-Stream output interface 96
    output m_axis_bram_96_tlast,
    output m_axis_bram_96_tvalid,
    output [C_OUTPUT_BRAM_96_DMWIDTH/8-1:0] m_axis_bram_96_tkeep,
    output [C_OUTPUT_BRAM_96_DMWIDTH/8-1:0] m_axis_bram_96_tstrb,
    output [C_OUTPUT_BRAM_96_DMWIDTH-1:0] m_axis_bram_96_tdata,
    input m_axis_bram_96_tready,
    input [C_OUTPUT_BRAM_96_ADDR_WIDTH-1:0] ap_bram_oarg_96_addr0,
    input [C_OUTPUT_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_din0,
    output [C_OUTPUT_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_dout0,
    input ap_bram_oarg_96_clk0,
    input ap_bram_oarg_96_rst0,
    input [C_OUTPUT_BRAM_96_WIDTH/8-1:0] ap_bram_oarg_96_we0,
    input ap_bram_oarg_96_en0,
    input [C_OUTPUT_BRAM_96_ADDR_WIDTH-1:0] ap_bram_oarg_96_addr1,
    input [C_OUTPUT_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_din1,
    output [C_OUTPUT_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_dout1,
    input ap_bram_oarg_96_clk1,
    input ap_bram_oarg_96_rst1,
    input [C_OUTPUT_BRAM_96_WIDTH/8-1:0] ap_bram_oarg_96_we1,
    input ap_bram_oarg_96_en1,
    //out AXI-Stream output interface 97
    output m_axis_bram_97_tlast,
    output m_axis_bram_97_tvalid,
    output [C_OUTPUT_BRAM_97_DMWIDTH/8-1:0] m_axis_bram_97_tkeep,
    output [C_OUTPUT_BRAM_97_DMWIDTH/8-1:0] m_axis_bram_97_tstrb,
    output [C_OUTPUT_BRAM_97_DMWIDTH-1:0] m_axis_bram_97_tdata,
    input m_axis_bram_97_tready,
    input [C_OUTPUT_BRAM_97_ADDR_WIDTH-1:0] ap_bram_oarg_97_addr0,
    input [C_OUTPUT_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_din0,
    output [C_OUTPUT_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_dout0,
    input ap_bram_oarg_97_clk0,
    input ap_bram_oarg_97_rst0,
    input [C_OUTPUT_BRAM_97_WIDTH/8-1:0] ap_bram_oarg_97_we0,
    input ap_bram_oarg_97_en0,
    input [C_OUTPUT_BRAM_97_ADDR_WIDTH-1:0] ap_bram_oarg_97_addr1,
    input [C_OUTPUT_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_din1,
    output [C_OUTPUT_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_dout1,
    input ap_bram_oarg_97_clk1,
    input ap_bram_oarg_97_rst1,
    input [C_OUTPUT_BRAM_97_WIDTH/8-1:0] ap_bram_oarg_97_we1,
    input ap_bram_oarg_97_en1,
    //out AXI-Stream output interface 98
    output m_axis_bram_98_tlast,
    output m_axis_bram_98_tvalid,
    output [C_OUTPUT_BRAM_98_DMWIDTH/8-1:0] m_axis_bram_98_tkeep,
    output [C_OUTPUT_BRAM_98_DMWIDTH/8-1:0] m_axis_bram_98_tstrb,
    output [C_OUTPUT_BRAM_98_DMWIDTH-1:0] m_axis_bram_98_tdata,
    input m_axis_bram_98_tready,
    input [C_OUTPUT_BRAM_98_ADDR_WIDTH-1:0] ap_bram_oarg_98_addr0,
    input [C_OUTPUT_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_din0,
    output [C_OUTPUT_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_dout0,
    input ap_bram_oarg_98_clk0,
    input ap_bram_oarg_98_rst0,
    input [C_OUTPUT_BRAM_98_WIDTH/8-1:0] ap_bram_oarg_98_we0,
    input ap_bram_oarg_98_en0,
    input [C_OUTPUT_BRAM_98_ADDR_WIDTH-1:0] ap_bram_oarg_98_addr1,
    input [C_OUTPUT_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_din1,
    output [C_OUTPUT_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_dout1,
    input ap_bram_oarg_98_clk1,
    input ap_bram_oarg_98_rst1,
    input [C_OUTPUT_BRAM_98_WIDTH/8-1:0] ap_bram_oarg_98_we1,
    input ap_bram_oarg_98_en1,
    //out AXI-Stream output interface 99
    output m_axis_bram_99_tlast,
    output m_axis_bram_99_tvalid,
    output [C_OUTPUT_BRAM_99_DMWIDTH/8-1:0] m_axis_bram_99_tkeep,
    output [C_OUTPUT_BRAM_99_DMWIDTH/8-1:0] m_axis_bram_99_tstrb,
    output [C_OUTPUT_BRAM_99_DMWIDTH-1:0] m_axis_bram_99_tdata,
    input m_axis_bram_99_tready,
    input [C_OUTPUT_BRAM_99_ADDR_WIDTH-1:0] ap_bram_oarg_99_addr0,
    input [C_OUTPUT_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_din0,
    output [C_OUTPUT_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_dout0,
    input ap_bram_oarg_99_clk0,
    input ap_bram_oarg_99_rst0,
    input [C_OUTPUT_BRAM_99_WIDTH/8-1:0] ap_bram_oarg_99_we0,
    input ap_bram_oarg_99_en0,
    input [C_OUTPUT_BRAM_99_ADDR_WIDTH-1:0] ap_bram_oarg_99_addr1,
    input [C_OUTPUT_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_din1,
    output [C_OUTPUT_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_dout1,
    input ap_bram_oarg_99_clk1,
    input ap_bram_oarg_99_rst1,
    input [C_OUTPUT_BRAM_99_WIDTH/8-1:0] ap_bram_oarg_99_we1,
    input ap_bram_oarg_99_en1,
    //out AXI-Stream output interface 100
    output m_axis_bram_100_tlast,
    output m_axis_bram_100_tvalid,
    output [C_OUTPUT_BRAM_100_DMWIDTH/8-1:0] m_axis_bram_100_tkeep,
    output [C_OUTPUT_BRAM_100_DMWIDTH/8-1:0] m_axis_bram_100_tstrb,
    output [C_OUTPUT_BRAM_100_DMWIDTH-1:0] m_axis_bram_100_tdata,
    input m_axis_bram_100_tready,
    input [C_OUTPUT_BRAM_100_ADDR_WIDTH-1:0] ap_bram_oarg_100_addr0,
    input [C_OUTPUT_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_din0,
    output [C_OUTPUT_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_dout0,
    input ap_bram_oarg_100_clk0,
    input ap_bram_oarg_100_rst0,
    input [C_OUTPUT_BRAM_100_WIDTH/8-1:0] ap_bram_oarg_100_we0,
    input ap_bram_oarg_100_en0,
    input [C_OUTPUT_BRAM_100_ADDR_WIDTH-1:0] ap_bram_oarg_100_addr1,
    input [C_OUTPUT_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_din1,
    output [C_OUTPUT_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_dout1,
    input ap_bram_oarg_100_clk1,
    input ap_bram_oarg_100_rst1,
    input [C_OUTPUT_BRAM_100_WIDTH/8-1:0] ap_bram_oarg_100_we1,
    input ap_bram_oarg_100_en1,
    //out AXI-Stream output interface 101
    output m_axis_bram_101_tlast,
    output m_axis_bram_101_tvalid,
    output [C_OUTPUT_BRAM_101_DMWIDTH/8-1:0] m_axis_bram_101_tkeep,
    output [C_OUTPUT_BRAM_101_DMWIDTH/8-1:0] m_axis_bram_101_tstrb,
    output [C_OUTPUT_BRAM_101_DMWIDTH-1:0] m_axis_bram_101_tdata,
    input m_axis_bram_101_tready,
    input [C_OUTPUT_BRAM_101_ADDR_WIDTH-1:0] ap_bram_oarg_101_addr0,
    input [C_OUTPUT_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_din0,
    output [C_OUTPUT_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_dout0,
    input ap_bram_oarg_101_clk0,
    input ap_bram_oarg_101_rst0,
    input [C_OUTPUT_BRAM_101_WIDTH/8-1:0] ap_bram_oarg_101_we0,
    input ap_bram_oarg_101_en0,
    input [C_OUTPUT_BRAM_101_ADDR_WIDTH-1:0] ap_bram_oarg_101_addr1,
    input [C_OUTPUT_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_din1,
    output [C_OUTPUT_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_dout1,
    input ap_bram_oarg_101_clk1,
    input ap_bram_oarg_101_rst1,
    input [C_OUTPUT_BRAM_101_WIDTH/8-1:0] ap_bram_oarg_101_we1,
    input ap_bram_oarg_101_en1,
    //out AXI-Stream output interface 102
    output m_axis_bram_102_tlast,
    output m_axis_bram_102_tvalid,
    output [C_OUTPUT_BRAM_102_DMWIDTH/8-1:0] m_axis_bram_102_tkeep,
    output [C_OUTPUT_BRAM_102_DMWIDTH/8-1:0] m_axis_bram_102_tstrb,
    output [C_OUTPUT_BRAM_102_DMWIDTH-1:0] m_axis_bram_102_tdata,
    input m_axis_bram_102_tready,
    input [C_OUTPUT_BRAM_102_ADDR_WIDTH-1:0] ap_bram_oarg_102_addr0,
    input [C_OUTPUT_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_din0,
    output [C_OUTPUT_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_dout0,
    input ap_bram_oarg_102_clk0,
    input ap_bram_oarg_102_rst0,
    input [C_OUTPUT_BRAM_102_WIDTH/8-1:0] ap_bram_oarg_102_we0,
    input ap_bram_oarg_102_en0,
    input [C_OUTPUT_BRAM_102_ADDR_WIDTH-1:0] ap_bram_oarg_102_addr1,
    input [C_OUTPUT_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_din1,
    output [C_OUTPUT_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_dout1,
    input ap_bram_oarg_102_clk1,
    input ap_bram_oarg_102_rst1,
    input [C_OUTPUT_BRAM_102_WIDTH/8-1:0] ap_bram_oarg_102_we1,
    input ap_bram_oarg_102_en1,
    //out AXI-Stream output interface 103
    output m_axis_bram_103_tlast,
    output m_axis_bram_103_tvalid,
    output [C_OUTPUT_BRAM_103_DMWIDTH/8-1:0] m_axis_bram_103_tkeep,
    output [C_OUTPUT_BRAM_103_DMWIDTH/8-1:0] m_axis_bram_103_tstrb,
    output [C_OUTPUT_BRAM_103_DMWIDTH-1:0] m_axis_bram_103_tdata,
    input m_axis_bram_103_tready,
    input [C_OUTPUT_BRAM_103_ADDR_WIDTH-1:0] ap_bram_oarg_103_addr0,
    input [C_OUTPUT_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_din0,
    output [C_OUTPUT_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_dout0,
    input ap_bram_oarg_103_clk0,
    input ap_bram_oarg_103_rst0,
    input [C_OUTPUT_BRAM_103_WIDTH/8-1:0] ap_bram_oarg_103_we0,
    input ap_bram_oarg_103_en0,
    input [C_OUTPUT_BRAM_103_ADDR_WIDTH-1:0] ap_bram_oarg_103_addr1,
    input [C_OUTPUT_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_din1,
    output [C_OUTPUT_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_dout1,
    input ap_bram_oarg_103_clk1,
    input ap_bram_oarg_103_rst1,
    input [C_OUTPUT_BRAM_103_WIDTH/8-1:0] ap_bram_oarg_103_we1,
    input ap_bram_oarg_103_en1,
    //out AXI-Stream output interface 104
    output m_axis_bram_104_tlast,
    output m_axis_bram_104_tvalid,
    output [C_OUTPUT_BRAM_104_DMWIDTH/8-1:0] m_axis_bram_104_tkeep,
    output [C_OUTPUT_BRAM_104_DMWIDTH/8-1:0] m_axis_bram_104_tstrb,
    output [C_OUTPUT_BRAM_104_DMWIDTH-1:0] m_axis_bram_104_tdata,
    input m_axis_bram_104_tready,
    input [C_OUTPUT_BRAM_104_ADDR_WIDTH-1:0] ap_bram_oarg_104_addr0,
    input [C_OUTPUT_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_din0,
    output [C_OUTPUT_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_dout0,
    input ap_bram_oarg_104_clk0,
    input ap_bram_oarg_104_rst0,
    input [C_OUTPUT_BRAM_104_WIDTH/8-1:0] ap_bram_oarg_104_we0,
    input ap_bram_oarg_104_en0,
    input [C_OUTPUT_BRAM_104_ADDR_WIDTH-1:0] ap_bram_oarg_104_addr1,
    input [C_OUTPUT_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_din1,
    output [C_OUTPUT_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_dout1,
    input ap_bram_oarg_104_clk1,
    input ap_bram_oarg_104_rst1,
    input [C_OUTPUT_BRAM_104_WIDTH/8-1:0] ap_bram_oarg_104_we1,
    input ap_bram_oarg_104_en1,
    //out AXI-Stream output interface 105
    output m_axis_bram_105_tlast,
    output m_axis_bram_105_tvalid,
    output [C_OUTPUT_BRAM_105_DMWIDTH/8-1:0] m_axis_bram_105_tkeep,
    output [C_OUTPUT_BRAM_105_DMWIDTH/8-1:0] m_axis_bram_105_tstrb,
    output [C_OUTPUT_BRAM_105_DMWIDTH-1:0] m_axis_bram_105_tdata,
    input m_axis_bram_105_tready,
    input [C_OUTPUT_BRAM_105_ADDR_WIDTH-1:0] ap_bram_oarg_105_addr0,
    input [C_OUTPUT_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_din0,
    output [C_OUTPUT_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_dout0,
    input ap_bram_oarg_105_clk0,
    input ap_bram_oarg_105_rst0,
    input [C_OUTPUT_BRAM_105_WIDTH/8-1:0] ap_bram_oarg_105_we0,
    input ap_bram_oarg_105_en0,
    input [C_OUTPUT_BRAM_105_ADDR_WIDTH-1:0] ap_bram_oarg_105_addr1,
    input [C_OUTPUT_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_din1,
    output [C_OUTPUT_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_dout1,
    input ap_bram_oarg_105_clk1,
    input ap_bram_oarg_105_rst1,
    input [C_OUTPUT_BRAM_105_WIDTH/8-1:0] ap_bram_oarg_105_we1,
    input ap_bram_oarg_105_en1,
    //out AXI-Stream output interface 106
    output m_axis_bram_106_tlast,
    output m_axis_bram_106_tvalid,
    output [C_OUTPUT_BRAM_106_DMWIDTH/8-1:0] m_axis_bram_106_tkeep,
    output [C_OUTPUT_BRAM_106_DMWIDTH/8-1:0] m_axis_bram_106_tstrb,
    output [C_OUTPUT_BRAM_106_DMWIDTH-1:0] m_axis_bram_106_tdata,
    input m_axis_bram_106_tready,
    input [C_OUTPUT_BRAM_106_ADDR_WIDTH-1:0] ap_bram_oarg_106_addr0,
    input [C_OUTPUT_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_din0,
    output [C_OUTPUT_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_dout0,
    input ap_bram_oarg_106_clk0,
    input ap_bram_oarg_106_rst0,
    input [C_OUTPUT_BRAM_106_WIDTH/8-1:0] ap_bram_oarg_106_we0,
    input ap_bram_oarg_106_en0,
    input [C_OUTPUT_BRAM_106_ADDR_WIDTH-1:0] ap_bram_oarg_106_addr1,
    input [C_OUTPUT_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_din1,
    output [C_OUTPUT_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_dout1,
    input ap_bram_oarg_106_clk1,
    input ap_bram_oarg_106_rst1,
    input [C_OUTPUT_BRAM_106_WIDTH/8-1:0] ap_bram_oarg_106_we1,
    input ap_bram_oarg_106_en1,
    //out AXI-Stream output interface 107
    output m_axis_bram_107_tlast,
    output m_axis_bram_107_tvalid,
    output [C_OUTPUT_BRAM_107_DMWIDTH/8-1:0] m_axis_bram_107_tkeep,
    output [C_OUTPUT_BRAM_107_DMWIDTH/8-1:0] m_axis_bram_107_tstrb,
    output [C_OUTPUT_BRAM_107_DMWIDTH-1:0] m_axis_bram_107_tdata,
    input m_axis_bram_107_tready,
    input [C_OUTPUT_BRAM_107_ADDR_WIDTH-1:0] ap_bram_oarg_107_addr0,
    input [C_OUTPUT_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_din0,
    output [C_OUTPUT_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_dout0,
    input ap_bram_oarg_107_clk0,
    input ap_bram_oarg_107_rst0,
    input [C_OUTPUT_BRAM_107_WIDTH/8-1:0] ap_bram_oarg_107_we0,
    input ap_bram_oarg_107_en0,
    input [C_OUTPUT_BRAM_107_ADDR_WIDTH-1:0] ap_bram_oarg_107_addr1,
    input [C_OUTPUT_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_din1,
    output [C_OUTPUT_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_dout1,
    input ap_bram_oarg_107_clk1,
    input ap_bram_oarg_107_rst1,
    input [C_OUTPUT_BRAM_107_WIDTH/8-1:0] ap_bram_oarg_107_we1,
    input ap_bram_oarg_107_en1,
    //out AXI-Stream output interface 108
    output m_axis_bram_108_tlast,
    output m_axis_bram_108_tvalid,
    output [C_OUTPUT_BRAM_108_DMWIDTH/8-1:0] m_axis_bram_108_tkeep,
    output [C_OUTPUT_BRAM_108_DMWIDTH/8-1:0] m_axis_bram_108_tstrb,
    output [C_OUTPUT_BRAM_108_DMWIDTH-1:0] m_axis_bram_108_tdata,
    input m_axis_bram_108_tready,
    input [C_OUTPUT_BRAM_108_ADDR_WIDTH-1:0] ap_bram_oarg_108_addr0,
    input [C_OUTPUT_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_din0,
    output [C_OUTPUT_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_dout0,
    input ap_bram_oarg_108_clk0,
    input ap_bram_oarg_108_rst0,
    input [C_OUTPUT_BRAM_108_WIDTH/8-1:0] ap_bram_oarg_108_we0,
    input ap_bram_oarg_108_en0,
    input [C_OUTPUT_BRAM_108_ADDR_WIDTH-1:0] ap_bram_oarg_108_addr1,
    input [C_OUTPUT_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_din1,
    output [C_OUTPUT_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_dout1,
    input ap_bram_oarg_108_clk1,
    input ap_bram_oarg_108_rst1,
    input [C_OUTPUT_BRAM_108_WIDTH/8-1:0] ap_bram_oarg_108_we1,
    input ap_bram_oarg_108_en1,
    //out AXI-Stream output interface 109
    output m_axis_bram_109_tlast,
    output m_axis_bram_109_tvalid,
    output [C_OUTPUT_BRAM_109_DMWIDTH/8-1:0] m_axis_bram_109_tkeep,
    output [C_OUTPUT_BRAM_109_DMWIDTH/8-1:0] m_axis_bram_109_tstrb,
    output [C_OUTPUT_BRAM_109_DMWIDTH-1:0] m_axis_bram_109_tdata,
    input m_axis_bram_109_tready,
    input [C_OUTPUT_BRAM_109_ADDR_WIDTH-1:0] ap_bram_oarg_109_addr0,
    input [C_OUTPUT_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_din0,
    output [C_OUTPUT_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_dout0,
    input ap_bram_oarg_109_clk0,
    input ap_bram_oarg_109_rst0,
    input [C_OUTPUT_BRAM_109_WIDTH/8-1:0] ap_bram_oarg_109_we0,
    input ap_bram_oarg_109_en0,
    input [C_OUTPUT_BRAM_109_ADDR_WIDTH-1:0] ap_bram_oarg_109_addr1,
    input [C_OUTPUT_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_din1,
    output [C_OUTPUT_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_dout1,
    input ap_bram_oarg_109_clk1,
    input ap_bram_oarg_109_rst1,
    input [C_OUTPUT_BRAM_109_WIDTH/8-1:0] ap_bram_oarg_109_we1,
    input ap_bram_oarg_109_en1,
    //out AXI-Stream output interface 110
    output m_axis_bram_110_tlast,
    output m_axis_bram_110_tvalid,
    output [C_OUTPUT_BRAM_110_DMWIDTH/8-1:0] m_axis_bram_110_tkeep,
    output [C_OUTPUT_BRAM_110_DMWIDTH/8-1:0] m_axis_bram_110_tstrb,
    output [C_OUTPUT_BRAM_110_DMWIDTH-1:0] m_axis_bram_110_tdata,
    input m_axis_bram_110_tready,
    input [C_OUTPUT_BRAM_110_ADDR_WIDTH-1:0] ap_bram_oarg_110_addr0,
    input [C_OUTPUT_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_din0,
    output [C_OUTPUT_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_dout0,
    input ap_bram_oarg_110_clk0,
    input ap_bram_oarg_110_rst0,
    input [C_OUTPUT_BRAM_110_WIDTH/8-1:0] ap_bram_oarg_110_we0,
    input ap_bram_oarg_110_en0,
    input [C_OUTPUT_BRAM_110_ADDR_WIDTH-1:0] ap_bram_oarg_110_addr1,
    input [C_OUTPUT_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_din1,
    output [C_OUTPUT_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_dout1,
    input ap_bram_oarg_110_clk1,
    input ap_bram_oarg_110_rst1,
    input [C_OUTPUT_BRAM_110_WIDTH/8-1:0] ap_bram_oarg_110_we1,
    input ap_bram_oarg_110_en1,
    //out AXI-Stream output interface 111
    output m_axis_bram_111_tlast,
    output m_axis_bram_111_tvalid,
    output [C_OUTPUT_BRAM_111_DMWIDTH/8-1:0] m_axis_bram_111_tkeep,
    output [C_OUTPUT_BRAM_111_DMWIDTH/8-1:0] m_axis_bram_111_tstrb,
    output [C_OUTPUT_BRAM_111_DMWIDTH-1:0] m_axis_bram_111_tdata,
    input m_axis_bram_111_tready,
    input [C_OUTPUT_BRAM_111_ADDR_WIDTH-1:0] ap_bram_oarg_111_addr0,
    input [C_OUTPUT_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_din0,
    output [C_OUTPUT_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_dout0,
    input ap_bram_oarg_111_clk0,
    input ap_bram_oarg_111_rst0,
    input [C_OUTPUT_BRAM_111_WIDTH/8-1:0] ap_bram_oarg_111_we0,
    input ap_bram_oarg_111_en0,
    input [C_OUTPUT_BRAM_111_ADDR_WIDTH-1:0] ap_bram_oarg_111_addr1,
    input [C_OUTPUT_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_din1,
    output [C_OUTPUT_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_dout1,
    input ap_bram_oarg_111_clk1,
    input ap_bram_oarg_111_rst1,
    input [C_OUTPUT_BRAM_111_WIDTH/8-1:0] ap_bram_oarg_111_we1,
    input ap_bram_oarg_111_en1,
    //out AXI-Stream output interface 112
    output m_axis_bram_112_tlast,
    output m_axis_bram_112_tvalid,
    output [C_OUTPUT_BRAM_112_DMWIDTH/8-1:0] m_axis_bram_112_tkeep,
    output [C_OUTPUT_BRAM_112_DMWIDTH/8-1:0] m_axis_bram_112_tstrb,
    output [C_OUTPUT_BRAM_112_DMWIDTH-1:0] m_axis_bram_112_tdata,
    input m_axis_bram_112_tready,
    input [C_OUTPUT_BRAM_112_ADDR_WIDTH-1:0] ap_bram_oarg_112_addr0,
    input [C_OUTPUT_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_din0,
    output [C_OUTPUT_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_dout0,
    input ap_bram_oarg_112_clk0,
    input ap_bram_oarg_112_rst0,
    input [C_OUTPUT_BRAM_112_WIDTH/8-1:0] ap_bram_oarg_112_we0,
    input ap_bram_oarg_112_en0,
    input [C_OUTPUT_BRAM_112_ADDR_WIDTH-1:0] ap_bram_oarg_112_addr1,
    input [C_OUTPUT_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_din1,
    output [C_OUTPUT_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_dout1,
    input ap_bram_oarg_112_clk1,
    input ap_bram_oarg_112_rst1,
    input [C_OUTPUT_BRAM_112_WIDTH/8-1:0] ap_bram_oarg_112_we1,
    input ap_bram_oarg_112_en1,
    //out AXI-Stream output interface 113
    output m_axis_bram_113_tlast,
    output m_axis_bram_113_tvalid,
    output [C_OUTPUT_BRAM_113_DMWIDTH/8-1:0] m_axis_bram_113_tkeep,
    output [C_OUTPUT_BRAM_113_DMWIDTH/8-1:0] m_axis_bram_113_tstrb,
    output [C_OUTPUT_BRAM_113_DMWIDTH-1:0] m_axis_bram_113_tdata,
    input m_axis_bram_113_tready,
    input [C_OUTPUT_BRAM_113_ADDR_WIDTH-1:0] ap_bram_oarg_113_addr0,
    input [C_OUTPUT_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_din0,
    output [C_OUTPUT_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_dout0,
    input ap_bram_oarg_113_clk0,
    input ap_bram_oarg_113_rst0,
    input [C_OUTPUT_BRAM_113_WIDTH/8-1:0] ap_bram_oarg_113_we0,
    input ap_bram_oarg_113_en0,
    input [C_OUTPUT_BRAM_113_ADDR_WIDTH-1:0] ap_bram_oarg_113_addr1,
    input [C_OUTPUT_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_din1,
    output [C_OUTPUT_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_dout1,
    input ap_bram_oarg_113_clk1,
    input ap_bram_oarg_113_rst1,
    input [C_OUTPUT_BRAM_113_WIDTH/8-1:0] ap_bram_oarg_113_we1,
    input ap_bram_oarg_113_en1,
    //out AXI-Stream output interface 114
    output m_axis_bram_114_tlast,
    output m_axis_bram_114_tvalid,
    output [C_OUTPUT_BRAM_114_DMWIDTH/8-1:0] m_axis_bram_114_tkeep,
    output [C_OUTPUT_BRAM_114_DMWIDTH/8-1:0] m_axis_bram_114_tstrb,
    output [C_OUTPUT_BRAM_114_DMWIDTH-1:0] m_axis_bram_114_tdata,
    input m_axis_bram_114_tready,
    input [C_OUTPUT_BRAM_114_ADDR_WIDTH-1:0] ap_bram_oarg_114_addr0,
    input [C_OUTPUT_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_din0,
    output [C_OUTPUT_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_dout0,
    input ap_bram_oarg_114_clk0,
    input ap_bram_oarg_114_rst0,
    input [C_OUTPUT_BRAM_114_WIDTH/8-1:0] ap_bram_oarg_114_we0,
    input ap_bram_oarg_114_en0,
    input [C_OUTPUT_BRAM_114_ADDR_WIDTH-1:0] ap_bram_oarg_114_addr1,
    input [C_OUTPUT_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_din1,
    output [C_OUTPUT_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_dout1,
    input ap_bram_oarg_114_clk1,
    input ap_bram_oarg_114_rst1,
    input [C_OUTPUT_BRAM_114_WIDTH/8-1:0] ap_bram_oarg_114_we1,
    input ap_bram_oarg_114_en1,
    //out AXI-Stream output interface 115
    output m_axis_bram_115_tlast,
    output m_axis_bram_115_tvalid,
    output [C_OUTPUT_BRAM_115_DMWIDTH/8-1:0] m_axis_bram_115_tkeep,
    output [C_OUTPUT_BRAM_115_DMWIDTH/8-1:0] m_axis_bram_115_tstrb,
    output [C_OUTPUT_BRAM_115_DMWIDTH-1:0] m_axis_bram_115_tdata,
    input m_axis_bram_115_tready,
    input [C_OUTPUT_BRAM_115_ADDR_WIDTH-1:0] ap_bram_oarg_115_addr0,
    input [C_OUTPUT_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_din0,
    output [C_OUTPUT_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_dout0,
    input ap_bram_oarg_115_clk0,
    input ap_bram_oarg_115_rst0,
    input [C_OUTPUT_BRAM_115_WIDTH/8-1:0] ap_bram_oarg_115_we0,
    input ap_bram_oarg_115_en0,
    input [C_OUTPUT_BRAM_115_ADDR_WIDTH-1:0] ap_bram_oarg_115_addr1,
    input [C_OUTPUT_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_din1,
    output [C_OUTPUT_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_dout1,
    input ap_bram_oarg_115_clk1,
    input ap_bram_oarg_115_rst1,
    input [C_OUTPUT_BRAM_115_WIDTH/8-1:0] ap_bram_oarg_115_we1,
    input ap_bram_oarg_115_en1,
    //out AXI-Stream output interface 116
    output m_axis_bram_116_tlast,
    output m_axis_bram_116_tvalid,
    output [C_OUTPUT_BRAM_116_DMWIDTH/8-1:0] m_axis_bram_116_tkeep,
    output [C_OUTPUT_BRAM_116_DMWIDTH/8-1:0] m_axis_bram_116_tstrb,
    output [C_OUTPUT_BRAM_116_DMWIDTH-1:0] m_axis_bram_116_tdata,
    input m_axis_bram_116_tready,
    input [C_OUTPUT_BRAM_116_ADDR_WIDTH-1:0] ap_bram_oarg_116_addr0,
    input [C_OUTPUT_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_din0,
    output [C_OUTPUT_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_dout0,
    input ap_bram_oarg_116_clk0,
    input ap_bram_oarg_116_rst0,
    input [C_OUTPUT_BRAM_116_WIDTH/8-1:0] ap_bram_oarg_116_we0,
    input ap_bram_oarg_116_en0,
    input [C_OUTPUT_BRAM_116_ADDR_WIDTH-1:0] ap_bram_oarg_116_addr1,
    input [C_OUTPUT_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_din1,
    output [C_OUTPUT_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_dout1,
    input ap_bram_oarg_116_clk1,
    input ap_bram_oarg_116_rst1,
    input [C_OUTPUT_BRAM_116_WIDTH/8-1:0] ap_bram_oarg_116_we1,
    input ap_bram_oarg_116_en1,
    //out AXI-Stream output interface 117
    output m_axis_bram_117_tlast,
    output m_axis_bram_117_tvalid,
    output [C_OUTPUT_BRAM_117_DMWIDTH/8-1:0] m_axis_bram_117_tkeep,
    output [C_OUTPUT_BRAM_117_DMWIDTH/8-1:0] m_axis_bram_117_tstrb,
    output [C_OUTPUT_BRAM_117_DMWIDTH-1:0] m_axis_bram_117_tdata,
    input m_axis_bram_117_tready,
    input [C_OUTPUT_BRAM_117_ADDR_WIDTH-1:0] ap_bram_oarg_117_addr0,
    input [C_OUTPUT_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_din0,
    output [C_OUTPUT_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_dout0,
    input ap_bram_oarg_117_clk0,
    input ap_bram_oarg_117_rst0,
    input [C_OUTPUT_BRAM_117_WIDTH/8-1:0] ap_bram_oarg_117_we0,
    input ap_bram_oarg_117_en0,
    input [C_OUTPUT_BRAM_117_ADDR_WIDTH-1:0] ap_bram_oarg_117_addr1,
    input [C_OUTPUT_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_din1,
    output [C_OUTPUT_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_dout1,
    input ap_bram_oarg_117_clk1,
    input ap_bram_oarg_117_rst1,
    input [C_OUTPUT_BRAM_117_WIDTH/8-1:0] ap_bram_oarg_117_we1,
    input ap_bram_oarg_117_en1,
    //out AXI-Stream output interface 118
    output m_axis_bram_118_tlast,
    output m_axis_bram_118_tvalid,
    output [C_OUTPUT_BRAM_118_DMWIDTH/8-1:0] m_axis_bram_118_tkeep,
    output [C_OUTPUT_BRAM_118_DMWIDTH/8-1:0] m_axis_bram_118_tstrb,
    output [C_OUTPUT_BRAM_118_DMWIDTH-1:0] m_axis_bram_118_tdata,
    input m_axis_bram_118_tready,
    input [C_OUTPUT_BRAM_118_ADDR_WIDTH-1:0] ap_bram_oarg_118_addr0,
    input [C_OUTPUT_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_din0,
    output [C_OUTPUT_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_dout0,
    input ap_bram_oarg_118_clk0,
    input ap_bram_oarg_118_rst0,
    input [C_OUTPUT_BRAM_118_WIDTH/8-1:0] ap_bram_oarg_118_we0,
    input ap_bram_oarg_118_en0,
    input [C_OUTPUT_BRAM_118_ADDR_WIDTH-1:0] ap_bram_oarg_118_addr1,
    input [C_OUTPUT_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_din1,
    output [C_OUTPUT_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_dout1,
    input ap_bram_oarg_118_clk1,
    input ap_bram_oarg_118_rst1,
    input [C_OUTPUT_BRAM_118_WIDTH/8-1:0] ap_bram_oarg_118_we1,
    input ap_bram_oarg_118_en1,
    //out AXI-Stream output interface 119
    output m_axis_bram_119_tlast,
    output m_axis_bram_119_tvalid,
    output [C_OUTPUT_BRAM_119_DMWIDTH/8-1:0] m_axis_bram_119_tkeep,
    output [C_OUTPUT_BRAM_119_DMWIDTH/8-1:0] m_axis_bram_119_tstrb,
    output [C_OUTPUT_BRAM_119_DMWIDTH-1:0] m_axis_bram_119_tdata,
    input m_axis_bram_119_tready,
    input [C_OUTPUT_BRAM_119_ADDR_WIDTH-1:0] ap_bram_oarg_119_addr0,
    input [C_OUTPUT_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_din0,
    output [C_OUTPUT_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_dout0,
    input ap_bram_oarg_119_clk0,
    input ap_bram_oarg_119_rst0,
    input [C_OUTPUT_BRAM_119_WIDTH/8-1:0] ap_bram_oarg_119_we0,
    input ap_bram_oarg_119_en0,
    input [C_OUTPUT_BRAM_119_ADDR_WIDTH-1:0] ap_bram_oarg_119_addr1,
    input [C_OUTPUT_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_din1,
    output [C_OUTPUT_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_dout1,
    input ap_bram_oarg_119_clk1,
    input ap_bram_oarg_119_rst1,
    input [C_OUTPUT_BRAM_119_WIDTH/8-1:0] ap_bram_oarg_119_we1,
    input ap_bram_oarg_119_en1,
    //out AXI-Stream output interface 120
    output m_axis_bram_120_tlast,
    output m_axis_bram_120_tvalid,
    output [C_OUTPUT_BRAM_120_DMWIDTH/8-1:0] m_axis_bram_120_tkeep,
    output [C_OUTPUT_BRAM_120_DMWIDTH/8-1:0] m_axis_bram_120_tstrb,
    output [C_OUTPUT_BRAM_120_DMWIDTH-1:0] m_axis_bram_120_tdata,
    input m_axis_bram_120_tready,
    input [C_OUTPUT_BRAM_120_ADDR_WIDTH-1:0] ap_bram_oarg_120_addr0,
    input [C_OUTPUT_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_din0,
    output [C_OUTPUT_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_dout0,
    input ap_bram_oarg_120_clk0,
    input ap_bram_oarg_120_rst0,
    input [C_OUTPUT_BRAM_120_WIDTH/8-1:0] ap_bram_oarg_120_we0,
    input ap_bram_oarg_120_en0,
    input [C_OUTPUT_BRAM_120_ADDR_WIDTH-1:0] ap_bram_oarg_120_addr1,
    input [C_OUTPUT_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_din1,
    output [C_OUTPUT_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_dout1,
    input ap_bram_oarg_120_clk1,
    input ap_bram_oarg_120_rst1,
    input [C_OUTPUT_BRAM_120_WIDTH/8-1:0] ap_bram_oarg_120_we1,
    input ap_bram_oarg_120_en1,
    //out AXI-Stream output interface 121
    output m_axis_bram_121_tlast,
    output m_axis_bram_121_tvalid,
    output [C_OUTPUT_BRAM_121_DMWIDTH/8-1:0] m_axis_bram_121_tkeep,
    output [C_OUTPUT_BRAM_121_DMWIDTH/8-1:0] m_axis_bram_121_tstrb,
    output [C_OUTPUT_BRAM_121_DMWIDTH-1:0] m_axis_bram_121_tdata,
    input m_axis_bram_121_tready,
    input [C_OUTPUT_BRAM_121_ADDR_WIDTH-1:0] ap_bram_oarg_121_addr0,
    input [C_OUTPUT_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_din0,
    output [C_OUTPUT_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_dout0,
    input ap_bram_oarg_121_clk0,
    input ap_bram_oarg_121_rst0,
    input [C_OUTPUT_BRAM_121_WIDTH/8-1:0] ap_bram_oarg_121_we0,
    input ap_bram_oarg_121_en0,
    input [C_OUTPUT_BRAM_121_ADDR_WIDTH-1:0] ap_bram_oarg_121_addr1,
    input [C_OUTPUT_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_din1,
    output [C_OUTPUT_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_dout1,
    input ap_bram_oarg_121_clk1,
    input ap_bram_oarg_121_rst1,
    input [C_OUTPUT_BRAM_121_WIDTH/8-1:0] ap_bram_oarg_121_we1,
    input ap_bram_oarg_121_en1,
    //out AXI-Stream output interface 122
    output m_axis_bram_122_tlast,
    output m_axis_bram_122_tvalid,
    output [C_OUTPUT_BRAM_122_DMWIDTH/8-1:0] m_axis_bram_122_tkeep,
    output [C_OUTPUT_BRAM_122_DMWIDTH/8-1:0] m_axis_bram_122_tstrb,
    output [C_OUTPUT_BRAM_122_DMWIDTH-1:0] m_axis_bram_122_tdata,
    input m_axis_bram_122_tready,
    input [C_OUTPUT_BRAM_122_ADDR_WIDTH-1:0] ap_bram_oarg_122_addr0,
    input [C_OUTPUT_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_din0,
    output [C_OUTPUT_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_dout0,
    input ap_bram_oarg_122_clk0,
    input ap_bram_oarg_122_rst0,
    input [C_OUTPUT_BRAM_122_WIDTH/8-1:0] ap_bram_oarg_122_we0,
    input ap_bram_oarg_122_en0,
    input [C_OUTPUT_BRAM_122_ADDR_WIDTH-1:0] ap_bram_oarg_122_addr1,
    input [C_OUTPUT_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_din1,
    output [C_OUTPUT_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_dout1,
    input ap_bram_oarg_122_clk1,
    input ap_bram_oarg_122_rst1,
    input [C_OUTPUT_BRAM_122_WIDTH/8-1:0] ap_bram_oarg_122_we1,
    input ap_bram_oarg_122_en1,
    //out AXI-Stream output interface 123
    output m_axis_bram_123_tlast,
    output m_axis_bram_123_tvalid,
    output [C_OUTPUT_BRAM_123_DMWIDTH/8-1:0] m_axis_bram_123_tkeep,
    output [C_OUTPUT_BRAM_123_DMWIDTH/8-1:0] m_axis_bram_123_tstrb,
    output [C_OUTPUT_BRAM_123_DMWIDTH-1:0] m_axis_bram_123_tdata,
    input m_axis_bram_123_tready,
    input [C_OUTPUT_BRAM_123_ADDR_WIDTH-1:0] ap_bram_oarg_123_addr0,
    input [C_OUTPUT_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_din0,
    output [C_OUTPUT_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_dout0,
    input ap_bram_oarg_123_clk0,
    input ap_bram_oarg_123_rst0,
    input [C_OUTPUT_BRAM_123_WIDTH/8-1:0] ap_bram_oarg_123_we0,
    input ap_bram_oarg_123_en0,
    input [C_OUTPUT_BRAM_123_ADDR_WIDTH-1:0] ap_bram_oarg_123_addr1,
    input [C_OUTPUT_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_din1,
    output [C_OUTPUT_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_dout1,
    input ap_bram_oarg_123_clk1,
    input ap_bram_oarg_123_rst1,
    input [C_OUTPUT_BRAM_123_WIDTH/8-1:0] ap_bram_oarg_123_we1,
    input ap_bram_oarg_123_en1,
    //out AXI-Stream output interface 124
    output m_axis_bram_124_tlast,
    output m_axis_bram_124_tvalid,
    output [C_OUTPUT_BRAM_124_DMWIDTH/8-1:0] m_axis_bram_124_tkeep,
    output [C_OUTPUT_BRAM_124_DMWIDTH/8-1:0] m_axis_bram_124_tstrb,
    output [C_OUTPUT_BRAM_124_DMWIDTH-1:0] m_axis_bram_124_tdata,
    input m_axis_bram_124_tready,
    input [C_OUTPUT_BRAM_124_ADDR_WIDTH-1:0] ap_bram_oarg_124_addr0,
    input [C_OUTPUT_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_din0,
    output [C_OUTPUT_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_dout0,
    input ap_bram_oarg_124_clk0,
    input ap_bram_oarg_124_rst0,
    input [C_OUTPUT_BRAM_124_WIDTH/8-1:0] ap_bram_oarg_124_we0,
    input ap_bram_oarg_124_en0,
    input [C_OUTPUT_BRAM_124_ADDR_WIDTH-1:0] ap_bram_oarg_124_addr1,
    input [C_OUTPUT_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_din1,
    output [C_OUTPUT_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_dout1,
    input ap_bram_oarg_124_clk1,
    input ap_bram_oarg_124_rst1,
    input [C_OUTPUT_BRAM_124_WIDTH/8-1:0] ap_bram_oarg_124_we1,
    input ap_bram_oarg_124_en1,
    //out AXI-Stream output interface 125
    output m_axis_bram_125_tlast,
    output m_axis_bram_125_tvalid,
    output [C_OUTPUT_BRAM_125_DMWIDTH/8-1:0] m_axis_bram_125_tkeep,
    output [C_OUTPUT_BRAM_125_DMWIDTH/8-1:0] m_axis_bram_125_tstrb,
    output [C_OUTPUT_BRAM_125_DMWIDTH-1:0] m_axis_bram_125_tdata,
    input m_axis_bram_125_tready,
    input [C_OUTPUT_BRAM_125_ADDR_WIDTH-1:0] ap_bram_oarg_125_addr0,
    input [C_OUTPUT_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_din0,
    output [C_OUTPUT_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_dout0,
    input ap_bram_oarg_125_clk0,
    input ap_bram_oarg_125_rst0,
    input [C_OUTPUT_BRAM_125_WIDTH/8-1:0] ap_bram_oarg_125_we0,
    input ap_bram_oarg_125_en0,
    input [C_OUTPUT_BRAM_125_ADDR_WIDTH-1:0] ap_bram_oarg_125_addr1,
    input [C_OUTPUT_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_din1,
    output [C_OUTPUT_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_dout1,
    input ap_bram_oarg_125_clk1,
    input ap_bram_oarg_125_rst1,
    input [C_OUTPUT_BRAM_125_WIDTH/8-1:0] ap_bram_oarg_125_we1,
    input ap_bram_oarg_125_en1,
    //out AXI-Stream output interface 126
    output m_axis_bram_126_tlast,
    output m_axis_bram_126_tvalid,
    output [C_OUTPUT_BRAM_126_DMWIDTH/8-1:0] m_axis_bram_126_tkeep,
    output [C_OUTPUT_BRAM_126_DMWIDTH/8-1:0] m_axis_bram_126_tstrb,
    output [C_OUTPUT_BRAM_126_DMWIDTH-1:0] m_axis_bram_126_tdata,
    input m_axis_bram_126_tready,
    input [C_OUTPUT_BRAM_126_ADDR_WIDTH-1:0] ap_bram_oarg_126_addr0,
    input [C_OUTPUT_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_din0,
    output [C_OUTPUT_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_dout0,
    input ap_bram_oarg_126_clk0,
    input ap_bram_oarg_126_rst0,
    input [C_OUTPUT_BRAM_126_WIDTH/8-1:0] ap_bram_oarg_126_we0,
    input ap_bram_oarg_126_en0,
    input [C_OUTPUT_BRAM_126_ADDR_WIDTH-1:0] ap_bram_oarg_126_addr1,
    input [C_OUTPUT_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_din1,
    output [C_OUTPUT_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_dout1,
    input ap_bram_oarg_126_clk1,
    input ap_bram_oarg_126_rst1,
    input [C_OUTPUT_BRAM_126_WIDTH/8-1:0] ap_bram_oarg_126_we1,
    input ap_bram_oarg_126_en1,
    //out AXI-Stream output interface 127
    output m_axis_bram_127_tlast,
    output m_axis_bram_127_tvalid,
    output [C_OUTPUT_BRAM_127_DMWIDTH/8-1:0] m_axis_bram_127_tkeep,
    output [C_OUTPUT_BRAM_127_DMWIDTH/8-1:0] m_axis_bram_127_tstrb,
    output [C_OUTPUT_BRAM_127_DMWIDTH-1:0] m_axis_bram_127_tdata,
    input m_axis_bram_127_tready,
    input [C_OUTPUT_BRAM_127_ADDR_WIDTH-1:0] ap_bram_oarg_127_addr0,
    input [C_OUTPUT_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_din0,
    output [C_OUTPUT_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_dout0,
    input ap_bram_oarg_127_clk0,
    input ap_bram_oarg_127_rst0,
    input [C_OUTPUT_BRAM_127_WIDTH/8-1:0] ap_bram_oarg_127_we0,
    input ap_bram_oarg_127_en0,
    input [C_OUTPUT_BRAM_127_ADDR_WIDTH-1:0] ap_bram_oarg_127_addr1,
    input [C_OUTPUT_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_din1,
    output [C_OUTPUT_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_dout1,
    input ap_bram_oarg_127_clk1,
    input ap_bram_oarg_127_rst1,
    input [C_OUTPUT_BRAM_127_WIDTH/8-1:0] ap_bram_oarg_127_we1,
    input ap_bram_oarg_127_en1
);

//adapter parameters
parameter C_ACC_RESET_POLARITY = 0;
parameter C_QUEUE_DEPTH = 16;

//scalar parameters
parameter C_N_INPUT_SCALARS = 0;
parameter C_N_OUTPUT_SCALARS = 0;
parameter C_FIFO_DEPTH = 16;
parameter C_HAS_RETURN = 0;
parameter [31:0] C_INPUT_SCALAR_0_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_1_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_2_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_3_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_4_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_5_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_6_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_7_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_8_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_9_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_10_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_11_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_12_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_13_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_14_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_15_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_16_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_17_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_18_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_19_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_20_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_21_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_22_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_23_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_24_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_25_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_26_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_27_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_28_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_29_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_30_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_31_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_32_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_33_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_34_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_35_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_36_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_37_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_38_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_39_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_40_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_41_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_42_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_43_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_44_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_45_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_46_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_47_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_48_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_49_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_50_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_51_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_52_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_53_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_54_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_55_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_56_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_57_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_58_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_59_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_60_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_61_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_62_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_63_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_64_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_65_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_66_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_67_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_68_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_69_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_70_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_71_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_72_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_73_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_74_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_75_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_76_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_77_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_78_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_79_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_80_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_81_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_82_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_83_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_84_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_85_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_86_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_87_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_88_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_89_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_90_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_91_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_92_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_93_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_94_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_95_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_96_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_97_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_98_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_99_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_100_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_101_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_102_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_103_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_104_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_105_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_106_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_107_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_108_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_109_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_110_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_111_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_112_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_113_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_114_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_115_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_116_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_117_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_118_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_119_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_120_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_121_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_122_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_123_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_124_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_125_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_126_WIDTH = 1;
parameter [31:0] C_INPUT_SCALAR_127_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_0_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_1_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_2_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_3_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_4_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_5_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_6_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_7_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_8_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_9_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_10_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_11_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_12_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_13_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_14_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_15_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_16_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_17_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_18_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_19_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_20_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_21_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_22_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_23_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_24_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_25_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_26_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_27_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_28_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_29_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_30_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_31_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_32_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_33_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_34_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_35_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_36_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_37_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_38_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_39_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_40_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_41_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_42_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_43_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_44_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_45_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_46_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_47_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_48_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_49_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_50_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_51_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_52_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_53_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_54_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_55_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_56_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_57_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_58_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_59_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_60_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_61_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_62_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_63_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_64_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_65_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_66_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_67_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_68_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_69_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_70_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_71_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_72_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_73_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_74_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_75_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_76_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_77_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_78_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_79_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_80_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_81_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_82_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_83_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_84_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_85_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_86_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_87_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_88_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_89_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_90_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_91_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_92_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_93_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_94_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_95_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_96_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_97_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_98_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_99_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_100_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_101_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_102_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_103_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_104_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_105_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_106_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_107_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_108_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_109_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_110_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_111_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_112_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_113_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_114_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_115_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_116_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_117_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_118_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_119_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_120_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_121_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_122_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_123_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_124_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_125_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_126_WIDTH = 1;
parameter [31:0]  C_OUTPUT_SCALAR_127_WIDTH = 1;

//fifo arg parameters
parameter C_NUM_INPUT_FIFOs = 0;                //number of input fifo interfaces on the accelerator
parameter C_NUM_OUTPUT_FIFOs = 0;               //number of output fifo interfaces on the accelerator
parameter [31:0] C_INPUT_FIFO_0_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_1_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_2_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_3_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_4_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_5_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_6_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_7_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_8_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_9_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_10_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_11_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_12_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_13_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_14_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_15_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_16_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_17_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_18_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_19_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_20_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_21_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_22_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_23_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_24_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_25_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_26_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_27_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_28_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_29_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_30_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_31_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_32_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_33_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_34_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_35_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_36_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_37_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_38_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_39_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_40_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_41_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_42_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_43_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_44_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_45_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_46_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_47_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_48_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_49_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_50_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_51_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_52_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_53_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_54_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_55_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_56_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_57_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_58_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_59_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_60_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_61_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_62_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_63_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_64_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_65_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_66_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_67_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_68_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_69_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_70_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_71_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_72_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_73_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_74_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_75_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_76_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_77_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_78_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_79_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_80_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_81_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_82_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_83_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_84_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_85_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_86_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_87_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_88_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_89_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_90_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_91_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_92_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_93_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_94_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_95_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_96_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_97_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_98_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_99_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_100_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_101_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_102_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_103_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_104_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_105_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_106_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_107_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_108_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_109_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_110_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_111_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_112_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_113_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_114_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_115_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_116_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_117_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_118_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_119_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_120_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_121_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_122_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_123_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_124_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_125_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_126_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_127_WIDTH = 8;     //width of input fifo interface on the accelerator
parameter [31:0] C_INPUT_FIFO_0_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_1_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_2_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_3_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_4_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_5_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_6_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_7_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_8_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_9_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_10_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_11_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_12_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_13_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_14_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_15_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_16_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_17_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_18_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_19_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_20_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_21_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_22_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_23_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_24_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_25_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_26_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_27_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_28_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_29_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_30_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_31_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_32_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_33_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_34_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_35_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_36_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_37_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_38_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_39_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_40_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_41_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_42_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_43_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_44_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_45_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_46_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_47_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_48_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_49_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_50_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_51_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_52_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_53_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_54_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_55_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_56_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_57_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_58_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_59_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_60_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_61_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_62_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_63_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_64_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_65_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_66_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_67_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_68_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_69_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_70_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_71_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_72_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_73_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_74_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_75_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_76_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_77_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_78_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_79_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_80_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_81_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_82_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_83_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_84_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_85_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_86_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_87_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_88_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_89_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_90_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_91_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_92_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_93_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_94_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_95_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_96_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_97_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_98_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_99_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_100_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_101_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_102_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_103_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_104_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_105_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_106_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_107_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_108_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_109_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_110_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_111_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_112_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_113_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_114_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_115_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_116_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_117_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_118_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_119_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_120_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_121_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_122_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_123_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_124_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_125_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_126_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_127_DEPTH = 16;      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_INPUT_FIFO_0_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_1_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_2_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_3_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_4_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_5_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_6_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_7_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_8_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_9_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_10_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_11_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_12_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_13_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_14_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_15_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_16_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_17_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_18_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_19_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_20_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_21_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_22_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_23_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_24_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_25_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_26_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_27_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_28_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_29_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_30_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_31_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_32_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_33_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_34_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_35_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_36_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_37_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_38_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_39_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_40_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_41_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_42_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_43_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_44_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_45_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_46_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_47_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_48_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_49_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_50_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_51_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_52_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_53_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_54_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_55_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_56_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_57_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_58_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_59_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_60_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_61_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_62_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_63_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_64_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_65_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_66_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_67_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_68_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_69_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_70_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_71_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_72_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_73_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_74_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_75_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_76_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_77_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_78_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_79_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_80_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_81_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_82_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_83_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_84_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_85_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_86_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_87_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_88_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_89_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_90_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_91_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_92_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_93_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_94_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_95_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_96_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_97_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_98_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_99_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_100_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_101_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_102_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_103_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_104_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_105_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_106_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_107_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_108_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_109_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_110_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_111_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_112_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_113_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_114_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_115_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_116_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_117_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_118_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_119_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_120_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_121_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_122_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_123_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_124_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_125_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_126_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_INPUT_FIFO_127_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input fifo interface
parameter [31:0] C_OUTPUT_FIFO_0_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_1_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_2_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_3_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_4_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_5_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_6_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_7_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_8_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_9_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_10_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_11_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_12_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_13_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_14_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_15_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_16_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_17_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_18_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_19_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_20_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_21_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_22_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_23_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_24_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_25_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_26_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_27_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_28_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_29_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_30_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_31_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_32_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_33_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_34_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_35_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_36_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_37_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_38_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_39_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_40_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_41_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_42_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_43_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_44_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_45_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_46_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_47_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_48_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_49_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_50_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_51_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_52_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_53_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_54_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_55_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_56_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_57_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_58_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_59_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_60_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_61_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_62_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_63_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_64_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_65_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_66_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_67_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_68_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_69_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_70_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_71_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_72_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_73_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_74_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_75_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_76_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_77_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_78_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_79_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_80_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_81_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_82_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_83_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_84_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_85_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_86_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_87_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_88_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_89_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_90_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_91_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_92_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_93_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_94_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_95_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_96_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_97_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_98_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_99_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_100_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_101_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_102_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_103_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_104_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_105_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_106_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_107_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_108_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_109_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_110_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_111_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_112_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_113_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_114_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_115_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_116_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_117_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_118_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_119_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_120_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_121_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_122_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_123_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_124_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_125_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_126_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_127_WIDTH = 8;    //width of output fifo interface on the accelerator
parameter [31:0] C_OUTPUT_FIFO_0_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_1_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_2_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_3_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_4_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_5_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_6_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_7_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_8_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_9_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_10_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_11_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_12_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_13_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_14_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_15_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_16_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_17_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_18_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_19_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_20_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_21_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_22_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_23_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_24_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_25_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_26_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_27_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_28_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_29_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_30_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_31_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_32_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_33_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_34_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_35_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_36_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_37_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_38_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_39_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_40_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_41_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_42_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_43_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_44_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_45_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_46_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_47_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_48_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_49_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_50_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_51_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_52_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_53_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_54_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_55_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_56_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_57_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_58_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_59_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_60_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_61_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_62_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_63_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_64_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_65_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_66_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_67_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_68_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_69_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_70_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_71_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_72_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_73_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_74_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_75_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_76_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_77_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_78_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_79_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_80_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_81_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_82_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_83_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_84_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_85_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_86_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_87_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_88_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_89_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_90_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_91_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_92_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_93_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_94_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_95_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_96_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_97_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_98_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_99_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_100_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_101_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_102_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_103_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_104_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_105_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_106_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_107_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_108_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_109_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_110_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_111_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_112_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_113_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_114_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_115_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_116_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_117_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_118_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_119_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_120_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_121_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_122_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_123_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_124_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_125_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_126_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_127_DEPTH = 16;     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
parameter [31:0] C_OUTPUT_FIFO_0_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_1_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_2_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_3_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_4_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_5_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_6_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_7_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_8_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_9_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_10_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_11_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_12_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_13_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_14_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_15_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_16_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_17_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_18_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_19_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_20_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_21_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_22_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_23_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_24_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_25_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_26_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_27_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_28_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_29_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_30_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_31_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_32_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_33_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_34_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_35_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_36_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_37_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_38_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_39_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_40_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_41_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_42_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_43_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_44_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_45_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_46_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_47_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_48_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_49_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_50_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_51_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_52_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_53_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_54_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_55_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_56_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_57_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_58_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_59_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_60_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_61_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_62_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_63_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_64_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_65_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_66_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_67_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_68_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_69_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_70_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_71_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_72_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_73_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_74_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_75_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_76_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_77_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_78_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_79_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_80_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_81_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_82_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_83_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_84_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_85_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_86_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_87_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_88_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_89_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_90_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_91_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_92_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_93_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_94_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_95_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_96_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_97_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_98_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_99_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_100_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_101_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_102_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_103_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_104_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_105_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_106_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_107_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_108_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_109_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_110_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_111_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_112_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_113_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_114_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_115_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_116_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_117_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_118_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_119_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_120_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_121_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_122_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_123_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_124_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_125_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_126_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface
parameter [31:0] C_OUTPUT_FIFO_127_DMWIDTH = 8;  //width of AXIS interface from DM to adapter for output fifo interface

//bram arg parameters
parameter C_NUM_INPUT_BRAMs = 0; 
parameter C_NUM_OUTPUT_BRAMs = 0; 
parameter C_INPUT_BRAM_0_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_1_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_2_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_3_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_4_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_5_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_6_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_7_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_8_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_9_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_10_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_11_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_12_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_13_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_14_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_15_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_16_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_17_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_18_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_19_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_20_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_21_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_22_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_23_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_24_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_25_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_26_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_27_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_28_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_29_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_30_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_31_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_32_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_33_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_34_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_35_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_36_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_37_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_38_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_39_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_40_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_41_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_42_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_43_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_44_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_45_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_46_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_47_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_48_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_49_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_50_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_51_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_52_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_53_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_54_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_55_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_56_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_57_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_58_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_59_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_60_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_61_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_62_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_63_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_64_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_65_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_66_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_67_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_68_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_69_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_70_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_71_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_72_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_73_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_74_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_75_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_76_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_77_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_78_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_79_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_80_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_81_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_82_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_83_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_84_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_85_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_86_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_87_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_88_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_89_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_90_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_91_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_92_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_93_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_94_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_95_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_96_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_97_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_98_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_99_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_100_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_101_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_102_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_103_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_104_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_105_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_106_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_107_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_108_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_109_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_110_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_111_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_112_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_113_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_114_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_115_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_116_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_117_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_118_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_119_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_120_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_121_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_122_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_123_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_124_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_125_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_126_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter C_INPUT_BRAM_127_PORTS = 1;            //number of bram ports (dual-ported, partitioned)
parameter [31:0] C_INPUT_BRAM_0_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_1_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_2_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_3_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_4_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_5_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_6_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_7_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_8_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_9_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_10_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_11_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_12_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_13_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_14_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_15_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_16_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_17_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_18_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_19_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_20_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_21_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_22_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_23_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_24_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_25_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_26_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_27_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_28_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_29_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_30_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_31_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_32_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_33_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_34_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_35_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_36_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_37_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_38_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_39_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_40_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_41_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_42_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_43_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_44_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_45_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_46_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_47_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_48_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_49_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_50_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_51_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_52_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_53_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_54_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_55_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_56_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_57_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_58_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_59_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_60_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_61_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_62_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_63_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_64_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_65_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_66_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_67_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_68_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_69_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_70_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_71_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_72_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_73_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_74_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_75_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_76_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_77_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_78_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_79_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_80_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_81_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_82_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_83_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_84_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_85_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_86_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_87_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_88_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_89_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_90_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_91_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_92_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_93_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_94_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_95_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_96_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_97_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_98_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_99_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_100_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_101_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_102_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_103_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_104_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_105_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_106_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_107_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_108_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_109_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_110_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_111_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_112_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_113_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_114_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_115_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_116_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_117_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_118_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_119_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_120_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_121_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_122_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_123_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_124_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_125_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_126_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_127_WIDTH = 8;     //width of input bram interface on the accelerator
parameter [31:0] C_INPUT_BRAM_0_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_1_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_2_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_3_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_4_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_5_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_6_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_7_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_8_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_9_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_10_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_11_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_12_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_13_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_14_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_15_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_16_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_17_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_18_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_19_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_20_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_21_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_22_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_23_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_24_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_25_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_26_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_27_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_28_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_29_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_30_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_31_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_32_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_33_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_34_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_35_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_36_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_37_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_38_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_39_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_40_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_41_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_42_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_43_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_44_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_45_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_46_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_47_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_48_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_49_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_50_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_51_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_52_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_53_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_54_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_55_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_56_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_57_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_58_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_59_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_60_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_61_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_62_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_63_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_64_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_65_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_66_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_67_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_68_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_69_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_70_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_71_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_72_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_73_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_74_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_75_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_76_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_77_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_78_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_79_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_80_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_81_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_82_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_83_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_84_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_85_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_86_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_87_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_88_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_89_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_90_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_91_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_92_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_93_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_94_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_95_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_96_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_97_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_98_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_99_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_100_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_101_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_102_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_103_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_104_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_105_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_106_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_107_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_108_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_109_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_110_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_111_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_112_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_113_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_114_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_115_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_116_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_117_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_118_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_119_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_120_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_121_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_122_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_123_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_124_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_125_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_126_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_127_DEPTH = 2;     //depth of BRAM in adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_0_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_1_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_2_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_3_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_4_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_5_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_6_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_7_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_8_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_9_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_10_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_11_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_12_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_13_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_14_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_15_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_16_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_17_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_18_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_19_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_20_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_21_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_22_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_23_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_24_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_25_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_26_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_27_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_28_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_29_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_30_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_31_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_32_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_33_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_34_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_35_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_36_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_37_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_38_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_39_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_40_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_41_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_42_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_43_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_44_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_45_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_46_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_47_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_48_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_49_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_50_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_51_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_52_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_53_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_54_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_55_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_56_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_57_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_58_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_59_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_60_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_61_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_62_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_63_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_64_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_65_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_66_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_67_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_68_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_69_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_70_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_71_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_72_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_73_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_74_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_75_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_76_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_77_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_78_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_79_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_80_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_81_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_82_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_83_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_84_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_85_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_86_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_87_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_88_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_89_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_90_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_91_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_92_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_93_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_94_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_95_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_96_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_97_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_98_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_99_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_100_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_101_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_102_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_103_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_104_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_105_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_106_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_107_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_108_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_109_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_110_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_111_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_112_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_113_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_114_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_115_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_116_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_117_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_118_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_119_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_120_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_121_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_122_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_123_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_124_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_125_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_126_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INPUT_BRAM_127_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for input bram interface
parameter [31:0] C_INOUT_BRAM_0_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_1_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_2_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_3_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_4_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_5_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_6_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_7_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_8_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_9_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_10_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_11_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_12_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_13_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_14_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_15_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_16_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_17_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_18_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_19_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_20_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_21_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_22_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_23_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_24_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_25_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_26_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_27_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_28_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_29_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_30_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_31_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_32_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_33_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_34_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_35_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_36_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_37_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_38_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_39_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_40_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_41_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_42_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_43_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_44_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_45_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_46_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_47_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_48_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_49_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_50_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_51_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_52_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_53_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_54_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_55_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_56_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_57_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_58_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_59_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_60_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_61_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_62_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_63_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_64_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_65_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_66_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_67_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_68_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_69_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_70_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_71_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_72_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_73_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_74_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_75_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_76_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_77_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_78_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_79_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_80_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_81_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_82_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_83_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_84_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_85_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_86_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_87_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_88_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_89_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_90_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_91_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_92_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_93_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_94_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_95_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_96_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_97_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_98_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_99_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_100_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_101_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_102_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_103_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_104_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_105_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_106_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_107_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_108_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_109_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_110_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_111_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_112_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_113_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_114_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_115_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_116_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_117_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_118_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_119_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_120_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_121_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_122_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_123_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_124_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_125_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_126_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [31:0] C_INOUT_BRAM_127_DMWIDTH = 8;   //width of AXIS interface from DM to adapter for inout (output) bram interface
parameter [0:0] C_BRAM_0_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_1_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_2_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_3_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_4_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_5_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_6_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_7_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_8_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_9_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_10_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_11_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_12_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_13_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_14_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_15_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_16_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_17_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_18_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_19_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_20_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_21_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_22_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_23_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_24_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_25_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_26_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_27_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_28_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_29_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_30_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_31_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_32_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_33_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_34_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_35_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_36_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_37_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_38_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_39_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_40_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_41_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_42_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_43_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_44_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_45_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_46_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_47_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_48_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_49_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_50_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_51_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_52_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_53_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_54_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_55_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_56_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_57_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_58_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_59_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_60_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_61_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_62_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_63_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_64_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_65_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_66_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_67_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_68_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_69_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_70_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_71_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_72_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_73_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_74_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_75_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_76_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_77_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_78_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_79_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_80_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_81_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_82_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_83_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_84_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_85_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_86_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_87_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_88_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_89_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_90_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_91_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_92_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_93_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_94_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_95_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_96_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_97_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_98_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_99_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_100_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_101_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_102_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_103_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_104_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_105_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_106_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_107_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_108_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_109_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_110_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_111_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_112_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_113_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_114_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_115_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_116_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_117_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_118_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_119_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_120_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_121_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_122_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_123_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_124_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_125_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_126_IS_INOUT = 0;         //enables the input bram also for output
parameter [0:0] C_BRAM_127_IS_INOUT = 0;         //enables the input bram also for output
parameter [31:0] C_INPUT_BRAM_0_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_1_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_2_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_3_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_4_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_5_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_6_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_7_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_8_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_9_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_10_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_11_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_12_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_13_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_14_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_15_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_16_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_17_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_18_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_19_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_20_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_21_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_22_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_23_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_24_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_25_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_26_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_27_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_28_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_29_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_30_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_31_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_32_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_33_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_34_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_35_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_36_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_37_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_38_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_39_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_40_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_41_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_42_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_43_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_44_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_45_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_46_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_47_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_48_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_49_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_50_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_51_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_52_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_53_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_54_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_55_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_56_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_57_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_58_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_59_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_60_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_61_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_62_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_63_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_64_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_65_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_66_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_67_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_68_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_69_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_70_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_71_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_72_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_73_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_74_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_75_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_76_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_77_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_78_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_79_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_80_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_81_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_82_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_83_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_84_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_85_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_86_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_87_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_88_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_89_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_90_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_91_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_92_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_93_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_94_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_95_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_96_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_97_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_98_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_99_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_100_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_101_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_102_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_103_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_104_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_105_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_106_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_107_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_108_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_109_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_110_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_111_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_112_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_113_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_114_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_115_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_116_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_117_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_118_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_119_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_120_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_121_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_122_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_123_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_124_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_125_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_126_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter [31:0] C_INPUT_BRAM_127_MB_DEPTH = 1;  //depth, number of copies of BRAM args
parameter C_OUTPUT_BRAM_0_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_1_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_2_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_3_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_4_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_5_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_6_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_7_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_8_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_9_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_10_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_11_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_12_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_13_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_14_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_15_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_16_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_17_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_18_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_19_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_20_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_21_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_22_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_23_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_24_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_25_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_26_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_27_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_28_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_29_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_30_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_31_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_32_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_33_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_34_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_35_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_36_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_37_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_38_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_39_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_40_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_41_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_42_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_43_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_44_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_45_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_46_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_47_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_48_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_49_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_50_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_51_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_52_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_53_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_54_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_55_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_56_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_57_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_58_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_59_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_60_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_61_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_62_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_63_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_64_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_65_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_66_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_67_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_68_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_69_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_70_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_71_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_72_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_73_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_74_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_75_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_76_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_77_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_78_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_79_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_80_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_81_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_82_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_83_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_84_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_85_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_86_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_87_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_88_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_89_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_90_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_91_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_92_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_93_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_94_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_95_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_96_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_97_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_98_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_99_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_100_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_101_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_102_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_103_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_104_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_105_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_106_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_107_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_108_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_109_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_110_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_111_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_112_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_113_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_114_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_115_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_116_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_117_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_118_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_119_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_120_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_121_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_122_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_123_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_124_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_125_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_126_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter C_OUTPUT_BRAM_127_PORTS = 1;           //number of bram ports (dual-ported, partitioned)
parameter [31:0] C_OUTPUT_BRAM_0_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_1_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_2_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_3_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_4_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_5_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_6_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_7_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_8_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_9_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_10_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_11_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_12_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_13_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_14_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_15_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_16_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_17_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_18_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_19_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_20_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_21_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_22_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_23_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_24_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_25_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_26_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_27_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_28_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_29_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_30_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_31_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_32_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_33_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_34_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_35_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_36_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_37_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_38_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_39_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_40_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_41_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_42_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_43_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_44_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_45_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_46_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_47_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_48_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_49_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_50_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_51_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_52_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_53_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_54_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_55_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_56_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_57_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_58_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_59_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_60_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_61_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_62_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_63_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_64_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_65_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_66_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_67_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_68_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_69_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_70_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_71_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_72_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_73_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_74_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_75_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_76_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_77_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_78_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_79_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_80_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_81_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_82_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_83_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_84_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_85_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_86_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_87_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_88_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_89_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_90_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_91_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_92_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_93_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_94_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_95_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_96_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_97_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_98_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_99_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_100_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_101_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_102_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_103_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_104_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_105_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_106_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_107_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_108_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_109_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_110_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_111_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_112_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_113_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_114_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_115_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_116_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_117_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_118_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_119_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_120_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_121_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_122_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_123_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_124_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_125_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_126_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_127_WIDTH = 8;    //width of output bram interface on the accelerator
parameter [31:0] C_OUTPUT_BRAM_0_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_1_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_2_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_3_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_4_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_5_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_6_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_7_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_8_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_9_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_10_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_11_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_12_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_13_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_14_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_15_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_16_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_17_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_18_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_19_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_20_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_21_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_22_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_23_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_24_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_25_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_26_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_27_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_28_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_29_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_30_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_31_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_32_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_33_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_34_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_35_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_36_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_37_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_38_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_39_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_40_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_41_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_42_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_43_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_44_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_45_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_46_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_47_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_48_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_49_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_50_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_51_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_52_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_53_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_54_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_55_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_56_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_57_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_58_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_59_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_60_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_61_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_62_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_63_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_64_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_65_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_66_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_67_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_68_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_69_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_70_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_71_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_72_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_73_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_74_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_75_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_76_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_77_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_78_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_79_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_80_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_81_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_82_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_83_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_84_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_85_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_86_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_87_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_88_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_89_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_90_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_91_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_92_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_93_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_94_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_95_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_96_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_97_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_98_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_99_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_100_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_101_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_102_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_103_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_104_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_105_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_106_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_107_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_108_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_109_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_110_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_111_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_112_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_113_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_114_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_115_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_116_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_117_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_118_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_119_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_120_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_121_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_122_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_123_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_124_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_125_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_126_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_127_DEPTH = 2;    //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_0_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_1_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_2_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_3_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_4_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_5_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_6_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_7_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_8_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_9_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_10_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_11_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_12_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_13_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_14_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_15_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_16_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_17_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_18_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_19_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_20_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_21_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_22_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_23_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_24_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_25_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_26_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_27_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_28_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_29_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_30_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_31_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_32_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_33_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_34_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_35_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_36_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_37_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_38_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_39_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_40_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_41_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_42_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_43_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_44_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_45_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_46_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_47_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_48_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_49_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_50_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_51_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_52_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_53_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_54_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_55_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_56_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_57_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_58_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_59_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_60_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_61_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_62_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_63_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_64_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_65_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_66_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_67_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_68_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_69_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_70_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_71_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_72_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_73_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_74_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_75_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_76_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_77_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_78_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_79_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_80_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_81_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_82_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_83_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_84_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_85_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_86_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_87_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_88_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_89_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_90_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_91_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_92_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_93_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_94_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_95_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_96_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_97_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_98_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_99_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_100_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_101_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_102_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_103_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_104_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_105_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_106_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_107_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_108_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_109_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_110_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_111_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_112_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_113_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_114_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_115_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_116_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_117_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_118_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_119_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_120_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_121_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_122_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_123_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_124_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_125_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_126_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_127_DMWIDTH = 8;  //width of AXIS interface from adapter to DM for output bram interface
parameter [31:0] C_OUTPUT_BRAM_0_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_1_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_2_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_3_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_4_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_5_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_6_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_7_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_8_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_9_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_10_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_11_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_12_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_13_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_14_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_15_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_16_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_17_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_18_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_19_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_20_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_21_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_22_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_23_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_24_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_25_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_26_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_27_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_28_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_29_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_30_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_31_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_32_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_33_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_34_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_35_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_36_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_37_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_38_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_39_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_40_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_41_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_42_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_43_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_44_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_45_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_46_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_47_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_48_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_49_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_50_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_51_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_52_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_53_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_54_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_55_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_56_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_57_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_58_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_59_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_60_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_61_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_62_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_63_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_64_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_65_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_66_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_67_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_68_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_69_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_70_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_71_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_72_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_73_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_74_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_75_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_76_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_77_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_78_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_79_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_80_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_81_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_82_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_83_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_84_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_85_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_86_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_87_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_88_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_89_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_90_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_91_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_92_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_93_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_94_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_95_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_96_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_97_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_98_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_99_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_100_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_101_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_102_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_103_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_104_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_105_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_106_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_107_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_108_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_109_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_110_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_111_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_112_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_113_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_114_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_115_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_116_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_117_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_118_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_119_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_120_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_121_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_122_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_123_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_124_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_125_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_126_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface
parameter [31:0] C_OUTPUT_BRAM_127_MB_DEPTH = 1; //depth of BRAM in adapter for output bram interface

parameter C_INPUT_BRAM_0_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_1_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_2_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_3_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_4_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_5_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_6_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_7_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_8_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_9_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_10_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_11_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_12_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_13_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_14_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_15_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_16_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_17_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_18_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_19_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_20_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_21_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_22_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_23_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_24_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_25_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_26_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_27_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_28_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_29_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_30_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_31_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_32_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_33_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_34_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_35_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_36_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_37_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_38_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_39_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_40_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_41_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_42_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_43_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_44_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_45_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_46_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_47_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_48_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_49_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_50_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_51_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_52_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_53_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_54_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_55_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_56_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_57_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_58_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_59_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_60_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_61_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_62_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_63_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_64_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_65_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_66_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_67_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_68_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_69_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_70_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_71_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_72_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_73_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_74_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_75_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_76_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_77_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_78_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_79_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_80_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_81_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_82_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_83_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_84_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_85_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_86_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_87_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_88_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_89_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_90_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_91_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_92_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_93_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_94_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_95_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_96_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_97_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_98_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_99_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_100_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_101_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_102_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_103_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_104_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_105_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_106_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_107_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_108_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_109_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_110_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_111_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_112_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_113_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_114_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_115_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_116_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_117_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_118_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_119_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_120_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_121_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_122_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_123_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_124_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_125_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_126_ADDR_WIDTH = 1;
parameter C_INPUT_BRAM_127_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_0_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_1_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_2_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_3_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_4_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_5_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_6_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_7_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_8_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_9_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_10_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_11_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_12_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_13_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_14_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_15_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_16_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_17_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_18_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_19_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_20_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_21_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_22_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_23_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_24_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_25_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_26_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_27_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_28_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_29_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_30_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_31_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_32_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_33_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_34_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_35_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_36_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_37_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_38_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_39_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_40_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_41_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_42_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_43_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_44_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_45_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_46_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_47_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_48_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_49_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_50_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_51_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_52_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_53_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_54_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_55_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_56_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_57_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_58_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_59_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_60_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_61_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_62_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_63_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_64_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_65_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_66_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_67_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_68_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_69_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_70_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_71_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_72_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_73_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_74_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_75_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_76_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_77_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_78_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_79_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_80_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_81_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_82_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_83_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_84_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_85_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_86_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_87_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_88_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_89_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_90_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_91_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_92_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_93_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_94_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_95_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_96_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_97_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_98_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_99_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_100_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_101_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_102_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_103_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_104_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_105_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_106_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_107_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_108_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_109_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_110_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_111_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_112_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_113_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_114_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_115_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_116_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_117_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_118_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_119_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_120_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_121_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_122_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_123_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_124_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_125_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_126_ADDR_WIDTH = 1;
parameter C_OUTPUT_BRAM_127_ADDR_WIDTH = 1;

    //scalar interface 
    wire [31:0] scalar_write_addr;
    wire [31:0] scalar_read_addr;
    wire [31:0] scalar_din;
    wire scalar_we;
    wire scalar_re;
    wire [31:0] scalar_dout;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_next;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_fifo_empty;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_fifo_full;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_fifo_empty;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_fifo_full;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_empty;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_dout;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_read;
    
    //wire in bram control interface
    wire inbram_ctrl_allow;
    wire [C_NUM_INPUT_BRAMs-1:0] inbram_ctrl_ready;
    wire [C_NUM_INPUT_BRAMs-1:0] inoutbram_ctrl_ready;
    wire [C_NUM_INPUT_BRAMs*32-1:0] inbram_depth;
    
    //wire in fifo control interface
    wire infifo_ctrl_allow;
    
    //wire out bram control interface
    wire outbram_ctrl_allow;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_ctrl_ready;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_ctrl_canstart;
    wire [C_NUM_OUTPUT_BRAMs*32-1:0] outbram_depth;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_depth_write;
    
    //wire out fifo control interface
    wire outfifo_ctrl_allow;

    adapter #(
        .C_ACC_RESET_POLARITY(C_ACC_RESET_POLARITY),
        .C_NUM_INPUT_SCALARS(C_N_INPUT_SCALARS),
        .C_NUM_OUTPUT_SCALARS(C_N_OUTPUT_SCALARS),
        .C_QUEUE_DEPTH(C_QUEUE_DEPTH),
        .C_NUM_INPUT_FIFOs(C_NUM_INPUT_FIFOs),
        .C_NUM_OUTPUT_FIFOs(C_NUM_OUTPUT_FIFOs),
        .C_NUM_INPUT_BRAMs(C_NUM_INPUT_BRAMs),
        .C_NUM_OUTPUT_BRAMs(C_NUM_OUTPUT_BRAMs)
    ) adapter_i (
        .S_AXI_ACLK(s_axi_aclk),
        .S_AXI_ARESETN(s_axi_aresetn),
        .S_AXI_AWADDR(S_AXI_AWADDR),
        .S_AXI_AWPROT(S_AXI_AWPROT),
        .S_AXI_AWVALID(S_AXI_AWVALID),
        .S_AXI_AWREADY(S_AXI_AWREADY),
        .S_AXI_WDATA(S_AXI_WDATA),
        .S_AXI_WSTRB(S_AXI_WSTRB),
        .S_AXI_WVALID(S_AXI_WVALID),
        .S_AXI_WREADY(S_AXI_WREADY),
        .S_AXI_BRESP(S_AXI_BRESP),
        .S_AXI_BVALID(S_AXI_BVALID),
        .S_AXI_BREADY(S_AXI_BREADY),
        .S_AXI_ARADDR(S_AXI_ARADDR),
        .S_AXI_ARPROT(S_AXI_ARPROT),
        .S_AXI_ARVALID(S_AXI_ARVALID),
        .S_AXI_ARREADY(S_AXI_ARREADY),
        .S_AXI_RDATA(S_AXI_RDATA),
        .S_AXI_RRESP(S_AXI_RRESP),
        .S_AXI_RVALID(S_AXI_RVALID),
        .S_AXI_RREADY(S_AXI_RREADY),
        .acc_clk(aclk),
        .acc_rstn(resetn),
        .ap_rst(aresetn),
        .ap_start(ap_start),
        .ap_start_single(ap_start_single),
        .ap_idle(ap_idle),
        .ap_done(ap_done),
        .ap_ready(ap_ready),
        .ap_continue(ap_continue),
        .ap_clk(ap_clk),
        .scalar_write_addr(scalar_write_addr),
        .scalar_read_addr(scalar_read_addr),
        .scalar_din(scalar_din),
        .scalar_we(scalar_we),
        .scalar_re(scalar_re),
        .scalar_dout(scalar_dout),
        .inscalar_next(inscalar_next),
        .inscalar_fifo_empty(inscalar_fifo_empty),
        .inscalar_fifo_full(inscalar_fifo_full),
        .outscalar_fifo_empty(outscalar_fifo_empty),
        .outscalar_fifo_full(outscalar_fifo_full),
        .outscalar_null_empty(outscalar_null_empty),
        .outscalar_null_dout(outscalar_null_dout),
        .outscalar_null_read(outscalar_null_read),
        .inbram_ctrl_allow(inbram_ctrl_allow),
        .inbram_ctrl_ready(inbram_ctrl_ready),
        .inoutbram_ctrl_ready(inoutbram_ctrl_ready),
        .infifo_ctrl_allow(infifo_ctrl_allow),
        .outbram_ctrl_allow(outbram_ctrl_allow),
        .outbram_ctrl_ready(outbram_ctrl_ready),
        .outbram_ctrl_canstart(outbram_ctrl_canstart),
        .outbram_depth(outbram_depth),
        .outbram_depth_write(outbram_depth_write),
        .outfifo_ctrl_allow(outfifo_ctrl_allow)
    );
    
    scalar #(
        .C_NUM_INSCALARS(C_N_INPUT_SCALARS),
        .C_NUM_OUTSCALARS(C_N_OUTPUT_SCALARS),
        .C_FIFO_DEPTH(C_FIFO_DEPTH),
        .C_HAS_RETURN(C_HAS_RETURN),
        .C_INSCALAR_0_BITS(C_INPUT_SCALAR_0_WIDTH),
        .C_INSCALAR_1_BITS(C_INPUT_SCALAR_1_WIDTH),
        .C_INSCALAR_2_BITS(C_INPUT_SCALAR_2_WIDTH),
        .C_INSCALAR_3_BITS(C_INPUT_SCALAR_3_WIDTH),
        .C_INSCALAR_4_BITS(C_INPUT_SCALAR_4_WIDTH),
        .C_INSCALAR_5_BITS(C_INPUT_SCALAR_5_WIDTH),
        .C_INSCALAR_6_BITS(C_INPUT_SCALAR_6_WIDTH),
        .C_INSCALAR_7_BITS(C_INPUT_SCALAR_7_WIDTH),
        .C_INSCALAR_8_BITS(C_INPUT_SCALAR_8_WIDTH),
        .C_INSCALAR_9_BITS(C_INPUT_SCALAR_9_WIDTH),
        .C_INSCALAR_10_BITS(C_INPUT_SCALAR_10_WIDTH),
        .C_INSCALAR_11_BITS(C_INPUT_SCALAR_11_WIDTH),
        .C_INSCALAR_12_BITS(C_INPUT_SCALAR_12_WIDTH),
        .C_INSCALAR_13_BITS(C_INPUT_SCALAR_13_WIDTH),
        .C_INSCALAR_14_BITS(C_INPUT_SCALAR_14_WIDTH),
        .C_INSCALAR_15_BITS(C_INPUT_SCALAR_15_WIDTH),
        .C_INSCALAR_16_BITS(C_INPUT_SCALAR_16_WIDTH),
        .C_INSCALAR_17_BITS(C_INPUT_SCALAR_17_WIDTH),
        .C_INSCALAR_18_BITS(C_INPUT_SCALAR_18_WIDTH),
        .C_INSCALAR_19_BITS(C_INPUT_SCALAR_19_WIDTH),
        .C_INSCALAR_20_BITS(C_INPUT_SCALAR_20_WIDTH),
        .C_INSCALAR_21_BITS(C_INPUT_SCALAR_21_WIDTH),
        .C_INSCALAR_22_BITS(C_INPUT_SCALAR_22_WIDTH),
        .C_INSCALAR_23_BITS(C_INPUT_SCALAR_23_WIDTH),
        .C_INSCALAR_24_BITS(C_INPUT_SCALAR_24_WIDTH),
        .C_INSCALAR_25_BITS(C_INPUT_SCALAR_25_WIDTH),
        .C_INSCALAR_26_BITS(C_INPUT_SCALAR_26_WIDTH),
        .C_INSCALAR_27_BITS(C_INPUT_SCALAR_27_WIDTH),
        .C_INSCALAR_28_BITS(C_INPUT_SCALAR_28_WIDTH),
        .C_INSCALAR_29_BITS(C_INPUT_SCALAR_29_WIDTH),
        .C_INSCALAR_30_BITS(C_INPUT_SCALAR_30_WIDTH),
        .C_INSCALAR_31_BITS(C_INPUT_SCALAR_31_WIDTH),
        .C_INSCALAR_32_BITS(C_INPUT_SCALAR_32_WIDTH),
        .C_INSCALAR_33_BITS(C_INPUT_SCALAR_33_WIDTH),
        .C_INSCALAR_34_BITS(C_INPUT_SCALAR_34_WIDTH),
        .C_INSCALAR_35_BITS(C_INPUT_SCALAR_35_WIDTH),
        .C_INSCALAR_36_BITS(C_INPUT_SCALAR_36_WIDTH),
        .C_INSCALAR_37_BITS(C_INPUT_SCALAR_37_WIDTH),
        .C_INSCALAR_38_BITS(C_INPUT_SCALAR_38_WIDTH),
        .C_INSCALAR_39_BITS(C_INPUT_SCALAR_39_WIDTH),
        .C_INSCALAR_40_BITS(C_INPUT_SCALAR_40_WIDTH),
        .C_INSCALAR_41_BITS(C_INPUT_SCALAR_41_WIDTH),
        .C_INSCALAR_42_BITS(C_INPUT_SCALAR_42_WIDTH),
        .C_INSCALAR_43_BITS(C_INPUT_SCALAR_43_WIDTH),
        .C_INSCALAR_44_BITS(C_INPUT_SCALAR_44_WIDTH),
        .C_INSCALAR_45_BITS(C_INPUT_SCALAR_45_WIDTH),
        .C_INSCALAR_46_BITS(C_INPUT_SCALAR_46_WIDTH),
        .C_INSCALAR_47_BITS(C_INPUT_SCALAR_47_WIDTH),
        .C_INSCALAR_48_BITS(C_INPUT_SCALAR_48_WIDTH),
        .C_INSCALAR_49_BITS(C_INPUT_SCALAR_49_WIDTH),
        .C_INSCALAR_50_BITS(C_INPUT_SCALAR_50_WIDTH),
        .C_INSCALAR_51_BITS(C_INPUT_SCALAR_51_WIDTH),
        .C_INSCALAR_52_BITS(C_INPUT_SCALAR_52_WIDTH),
        .C_INSCALAR_53_BITS(C_INPUT_SCALAR_53_WIDTH),
        .C_INSCALAR_54_BITS(C_INPUT_SCALAR_54_WIDTH),
        .C_INSCALAR_55_BITS(C_INPUT_SCALAR_55_WIDTH),
        .C_INSCALAR_56_BITS(C_INPUT_SCALAR_56_WIDTH),
        .C_INSCALAR_57_BITS(C_INPUT_SCALAR_57_WIDTH),
        .C_INSCALAR_58_BITS(C_INPUT_SCALAR_58_WIDTH),
        .C_INSCALAR_59_BITS(C_INPUT_SCALAR_59_WIDTH),
        .C_INSCALAR_60_BITS(C_INPUT_SCALAR_60_WIDTH),
        .C_INSCALAR_61_BITS(C_INPUT_SCALAR_61_WIDTH),
        .C_INSCALAR_62_BITS(C_INPUT_SCALAR_62_WIDTH),
        .C_INSCALAR_63_BITS(C_INPUT_SCALAR_63_WIDTH),
        .C_INSCALAR_64_BITS(C_INPUT_SCALAR_64_WIDTH),
        .C_INSCALAR_65_BITS(C_INPUT_SCALAR_65_WIDTH),
        .C_INSCALAR_66_BITS(C_INPUT_SCALAR_66_WIDTH),
        .C_INSCALAR_67_BITS(C_INPUT_SCALAR_67_WIDTH),
        .C_INSCALAR_68_BITS(C_INPUT_SCALAR_68_WIDTH),
        .C_INSCALAR_69_BITS(C_INPUT_SCALAR_69_WIDTH),
        .C_INSCALAR_70_BITS(C_INPUT_SCALAR_70_WIDTH),
        .C_INSCALAR_71_BITS(C_INPUT_SCALAR_71_WIDTH),
        .C_INSCALAR_72_BITS(C_INPUT_SCALAR_72_WIDTH),
        .C_INSCALAR_73_BITS(C_INPUT_SCALAR_73_WIDTH),
        .C_INSCALAR_74_BITS(C_INPUT_SCALAR_74_WIDTH),
        .C_INSCALAR_75_BITS(C_INPUT_SCALAR_75_WIDTH),
        .C_INSCALAR_76_BITS(C_INPUT_SCALAR_76_WIDTH),
        .C_INSCALAR_77_BITS(C_INPUT_SCALAR_77_WIDTH),
        .C_INSCALAR_78_BITS(C_INPUT_SCALAR_78_WIDTH),
        .C_INSCALAR_79_BITS(C_INPUT_SCALAR_79_WIDTH),
        .C_INSCALAR_80_BITS(C_INPUT_SCALAR_80_WIDTH),
        .C_INSCALAR_81_BITS(C_INPUT_SCALAR_81_WIDTH),
        .C_INSCALAR_82_BITS(C_INPUT_SCALAR_82_WIDTH),
        .C_INSCALAR_83_BITS(C_INPUT_SCALAR_83_WIDTH),
        .C_INSCALAR_84_BITS(C_INPUT_SCALAR_84_WIDTH),
        .C_INSCALAR_85_BITS(C_INPUT_SCALAR_85_WIDTH),
        .C_INSCALAR_86_BITS(C_INPUT_SCALAR_86_WIDTH),
        .C_INSCALAR_87_BITS(C_INPUT_SCALAR_87_WIDTH),
        .C_INSCALAR_88_BITS(C_INPUT_SCALAR_88_WIDTH),
        .C_INSCALAR_89_BITS(C_INPUT_SCALAR_89_WIDTH),
        .C_INSCALAR_90_BITS(C_INPUT_SCALAR_90_WIDTH),
        .C_INSCALAR_91_BITS(C_INPUT_SCALAR_91_WIDTH),
        .C_INSCALAR_92_BITS(C_INPUT_SCALAR_92_WIDTH),
        .C_INSCALAR_93_BITS(C_INPUT_SCALAR_93_WIDTH),
        .C_INSCALAR_94_BITS(C_INPUT_SCALAR_94_WIDTH),
        .C_INSCALAR_95_BITS(C_INPUT_SCALAR_95_WIDTH),
        .C_INSCALAR_96_BITS(C_INPUT_SCALAR_96_WIDTH),
        .C_INSCALAR_97_BITS(C_INPUT_SCALAR_97_WIDTH),
        .C_INSCALAR_98_BITS(C_INPUT_SCALAR_98_WIDTH),
        .C_INSCALAR_99_BITS(C_INPUT_SCALAR_99_WIDTH),
        .C_INSCALAR_100_BITS(C_INPUT_SCALAR_100_WIDTH),
        .C_INSCALAR_101_BITS(C_INPUT_SCALAR_101_WIDTH),
        .C_INSCALAR_102_BITS(C_INPUT_SCALAR_102_WIDTH),
        .C_INSCALAR_103_BITS(C_INPUT_SCALAR_103_WIDTH),
        .C_INSCALAR_104_BITS(C_INPUT_SCALAR_104_WIDTH),
        .C_INSCALAR_105_BITS(C_INPUT_SCALAR_105_WIDTH),
        .C_INSCALAR_106_BITS(C_INPUT_SCALAR_106_WIDTH),
        .C_INSCALAR_107_BITS(C_INPUT_SCALAR_107_WIDTH),
        .C_INSCALAR_108_BITS(C_INPUT_SCALAR_108_WIDTH),
        .C_INSCALAR_109_BITS(C_INPUT_SCALAR_109_WIDTH),
        .C_INSCALAR_110_BITS(C_INPUT_SCALAR_110_WIDTH),
        .C_INSCALAR_111_BITS(C_INPUT_SCALAR_111_WIDTH),
        .C_INSCALAR_112_BITS(C_INPUT_SCALAR_112_WIDTH),
        .C_INSCALAR_113_BITS(C_INPUT_SCALAR_113_WIDTH),
        .C_INSCALAR_114_BITS(C_INPUT_SCALAR_114_WIDTH),
        .C_INSCALAR_115_BITS(C_INPUT_SCALAR_115_WIDTH),
        .C_INSCALAR_116_BITS(C_INPUT_SCALAR_116_WIDTH),
        .C_INSCALAR_117_BITS(C_INPUT_SCALAR_117_WIDTH),
        .C_INSCALAR_118_BITS(C_INPUT_SCALAR_118_WIDTH),
        .C_INSCALAR_119_BITS(C_INPUT_SCALAR_119_WIDTH),
        .C_INSCALAR_120_BITS(C_INPUT_SCALAR_120_WIDTH),
        .C_INSCALAR_121_BITS(C_INPUT_SCALAR_121_WIDTH),
        .C_INSCALAR_122_BITS(C_INPUT_SCALAR_122_WIDTH),
        .C_INSCALAR_123_BITS(C_INPUT_SCALAR_123_WIDTH),
        .C_INSCALAR_124_BITS(C_INPUT_SCALAR_124_WIDTH),
        .C_INSCALAR_125_BITS(C_INPUT_SCALAR_125_WIDTH),
        .C_INSCALAR_126_BITS(C_INPUT_SCALAR_126_WIDTH),
        .C_INSCALAR_127_BITS(C_INPUT_SCALAR_127_WIDTH),
        .C_OUTSCALAR_0_BITS(C_OUTPUT_SCALAR_0_WIDTH),
        .C_OUTSCALAR_1_BITS(C_OUTPUT_SCALAR_1_WIDTH),
        .C_OUTSCALAR_2_BITS(C_OUTPUT_SCALAR_2_WIDTH),
        .C_OUTSCALAR_3_BITS(C_OUTPUT_SCALAR_3_WIDTH),
        .C_OUTSCALAR_4_BITS(C_OUTPUT_SCALAR_4_WIDTH),
        .C_OUTSCALAR_5_BITS(C_OUTPUT_SCALAR_5_WIDTH),
        .C_OUTSCALAR_6_BITS(C_OUTPUT_SCALAR_6_WIDTH),
        .C_OUTSCALAR_7_BITS(C_OUTPUT_SCALAR_7_WIDTH),
        .C_OUTSCALAR_8_BITS(C_OUTPUT_SCALAR_8_WIDTH),
        .C_OUTSCALAR_9_BITS(C_OUTPUT_SCALAR_9_WIDTH),
        .C_OUTSCALAR_10_BITS(C_OUTPUT_SCALAR_10_WIDTH),
        .C_OUTSCALAR_11_BITS(C_OUTPUT_SCALAR_11_WIDTH),
        .C_OUTSCALAR_12_BITS(C_OUTPUT_SCALAR_12_WIDTH),
        .C_OUTSCALAR_13_BITS(C_OUTPUT_SCALAR_13_WIDTH),
        .C_OUTSCALAR_14_BITS(C_OUTPUT_SCALAR_14_WIDTH),
        .C_OUTSCALAR_15_BITS(C_OUTPUT_SCALAR_15_WIDTH),
        .C_OUTSCALAR_16_BITS(C_OUTPUT_SCALAR_16_WIDTH),
        .C_OUTSCALAR_17_BITS(C_OUTPUT_SCALAR_17_WIDTH),
        .C_OUTSCALAR_18_BITS(C_OUTPUT_SCALAR_18_WIDTH),
        .C_OUTSCALAR_19_BITS(C_OUTPUT_SCALAR_19_WIDTH),
        .C_OUTSCALAR_20_BITS(C_OUTPUT_SCALAR_20_WIDTH),
        .C_OUTSCALAR_21_BITS(C_OUTPUT_SCALAR_21_WIDTH),
        .C_OUTSCALAR_22_BITS(C_OUTPUT_SCALAR_22_WIDTH),
        .C_OUTSCALAR_23_BITS(C_OUTPUT_SCALAR_23_WIDTH),
        .C_OUTSCALAR_24_BITS(C_OUTPUT_SCALAR_24_WIDTH),
        .C_OUTSCALAR_25_BITS(C_OUTPUT_SCALAR_25_WIDTH),
        .C_OUTSCALAR_26_BITS(C_OUTPUT_SCALAR_26_WIDTH),
        .C_OUTSCALAR_27_BITS(C_OUTPUT_SCALAR_27_WIDTH),
        .C_OUTSCALAR_28_BITS(C_OUTPUT_SCALAR_28_WIDTH),
        .C_OUTSCALAR_29_BITS(C_OUTPUT_SCALAR_29_WIDTH),
        .C_OUTSCALAR_30_BITS(C_OUTPUT_SCALAR_30_WIDTH),
        .C_OUTSCALAR_31_BITS(C_OUTPUT_SCALAR_31_WIDTH),
        .C_OUTSCALAR_32_BITS(C_OUTPUT_SCALAR_32_WIDTH),
        .C_OUTSCALAR_33_BITS(C_OUTPUT_SCALAR_33_WIDTH),
        .C_OUTSCALAR_34_BITS(C_OUTPUT_SCALAR_34_WIDTH),
        .C_OUTSCALAR_35_BITS(C_OUTPUT_SCALAR_35_WIDTH),
        .C_OUTSCALAR_36_BITS(C_OUTPUT_SCALAR_36_WIDTH),
        .C_OUTSCALAR_37_BITS(C_OUTPUT_SCALAR_37_WIDTH),
        .C_OUTSCALAR_38_BITS(C_OUTPUT_SCALAR_38_WIDTH),
        .C_OUTSCALAR_39_BITS(C_OUTPUT_SCALAR_39_WIDTH),
        .C_OUTSCALAR_40_BITS(C_OUTPUT_SCALAR_40_WIDTH),
        .C_OUTSCALAR_41_BITS(C_OUTPUT_SCALAR_41_WIDTH),
        .C_OUTSCALAR_42_BITS(C_OUTPUT_SCALAR_42_WIDTH),
        .C_OUTSCALAR_43_BITS(C_OUTPUT_SCALAR_43_WIDTH),
        .C_OUTSCALAR_44_BITS(C_OUTPUT_SCALAR_44_WIDTH),
        .C_OUTSCALAR_45_BITS(C_OUTPUT_SCALAR_45_WIDTH),
        .C_OUTSCALAR_46_BITS(C_OUTPUT_SCALAR_46_WIDTH),
        .C_OUTSCALAR_47_BITS(C_OUTPUT_SCALAR_47_WIDTH),
        .C_OUTSCALAR_48_BITS(C_OUTPUT_SCALAR_48_WIDTH),
        .C_OUTSCALAR_49_BITS(C_OUTPUT_SCALAR_49_WIDTH),
        .C_OUTSCALAR_50_BITS(C_OUTPUT_SCALAR_50_WIDTH),
        .C_OUTSCALAR_51_BITS(C_OUTPUT_SCALAR_51_WIDTH),
        .C_OUTSCALAR_52_BITS(C_OUTPUT_SCALAR_52_WIDTH),
        .C_OUTSCALAR_53_BITS(C_OUTPUT_SCALAR_53_WIDTH),
        .C_OUTSCALAR_54_BITS(C_OUTPUT_SCALAR_54_WIDTH),
        .C_OUTSCALAR_55_BITS(C_OUTPUT_SCALAR_55_WIDTH),
        .C_OUTSCALAR_56_BITS(C_OUTPUT_SCALAR_56_WIDTH),
        .C_OUTSCALAR_57_BITS(C_OUTPUT_SCALAR_57_WIDTH),
        .C_OUTSCALAR_58_BITS(C_OUTPUT_SCALAR_58_WIDTH),
        .C_OUTSCALAR_59_BITS(C_OUTPUT_SCALAR_59_WIDTH),
        .C_OUTSCALAR_60_BITS(C_OUTPUT_SCALAR_60_WIDTH),
        .C_OUTSCALAR_61_BITS(C_OUTPUT_SCALAR_61_WIDTH),
        .C_OUTSCALAR_62_BITS(C_OUTPUT_SCALAR_62_WIDTH),
        .C_OUTSCALAR_63_BITS(C_OUTPUT_SCALAR_63_WIDTH),
        .C_OUTSCALAR_64_BITS(C_OUTPUT_SCALAR_64_WIDTH),
        .C_OUTSCALAR_65_BITS(C_OUTPUT_SCALAR_65_WIDTH),
        .C_OUTSCALAR_66_BITS(C_OUTPUT_SCALAR_66_WIDTH),
        .C_OUTSCALAR_67_BITS(C_OUTPUT_SCALAR_67_WIDTH),
        .C_OUTSCALAR_68_BITS(C_OUTPUT_SCALAR_68_WIDTH),
        .C_OUTSCALAR_69_BITS(C_OUTPUT_SCALAR_69_WIDTH),
        .C_OUTSCALAR_70_BITS(C_OUTPUT_SCALAR_70_WIDTH),
        .C_OUTSCALAR_71_BITS(C_OUTPUT_SCALAR_71_WIDTH),
        .C_OUTSCALAR_72_BITS(C_OUTPUT_SCALAR_72_WIDTH),
        .C_OUTSCALAR_73_BITS(C_OUTPUT_SCALAR_73_WIDTH),
        .C_OUTSCALAR_74_BITS(C_OUTPUT_SCALAR_74_WIDTH),
        .C_OUTSCALAR_75_BITS(C_OUTPUT_SCALAR_75_WIDTH),
        .C_OUTSCALAR_76_BITS(C_OUTPUT_SCALAR_76_WIDTH),
        .C_OUTSCALAR_77_BITS(C_OUTPUT_SCALAR_77_WIDTH),
        .C_OUTSCALAR_78_BITS(C_OUTPUT_SCALAR_78_WIDTH),
        .C_OUTSCALAR_79_BITS(C_OUTPUT_SCALAR_79_WIDTH),
        .C_OUTSCALAR_80_BITS(C_OUTPUT_SCALAR_80_WIDTH),
        .C_OUTSCALAR_81_BITS(C_OUTPUT_SCALAR_81_WIDTH),
        .C_OUTSCALAR_82_BITS(C_OUTPUT_SCALAR_82_WIDTH),
        .C_OUTSCALAR_83_BITS(C_OUTPUT_SCALAR_83_WIDTH),
        .C_OUTSCALAR_84_BITS(C_OUTPUT_SCALAR_84_WIDTH),
        .C_OUTSCALAR_85_BITS(C_OUTPUT_SCALAR_85_WIDTH),
        .C_OUTSCALAR_86_BITS(C_OUTPUT_SCALAR_86_WIDTH),
        .C_OUTSCALAR_87_BITS(C_OUTPUT_SCALAR_87_WIDTH),
        .C_OUTSCALAR_88_BITS(C_OUTPUT_SCALAR_88_WIDTH),
        .C_OUTSCALAR_89_BITS(C_OUTPUT_SCALAR_89_WIDTH),
        .C_OUTSCALAR_90_BITS(C_OUTPUT_SCALAR_90_WIDTH),
        .C_OUTSCALAR_91_BITS(C_OUTPUT_SCALAR_91_WIDTH),
        .C_OUTSCALAR_92_BITS(C_OUTPUT_SCALAR_92_WIDTH),
        .C_OUTSCALAR_93_BITS(C_OUTPUT_SCALAR_93_WIDTH),
        .C_OUTSCALAR_94_BITS(C_OUTPUT_SCALAR_94_WIDTH),
        .C_OUTSCALAR_95_BITS(C_OUTPUT_SCALAR_95_WIDTH),
        .C_OUTSCALAR_96_BITS(C_OUTPUT_SCALAR_96_WIDTH),
        .C_OUTSCALAR_97_BITS(C_OUTPUT_SCALAR_97_WIDTH),
        .C_OUTSCALAR_98_BITS(C_OUTPUT_SCALAR_98_WIDTH),
        .C_OUTSCALAR_99_BITS(C_OUTPUT_SCALAR_99_WIDTH),
        .C_OUTSCALAR_100_BITS(C_OUTPUT_SCALAR_100_WIDTH),
        .C_OUTSCALAR_101_BITS(C_OUTPUT_SCALAR_101_WIDTH),
        .C_OUTSCALAR_102_BITS(C_OUTPUT_SCALAR_102_WIDTH),
        .C_OUTSCALAR_103_BITS(C_OUTPUT_SCALAR_103_WIDTH),
        .C_OUTSCALAR_104_BITS(C_OUTPUT_SCALAR_104_WIDTH),
        .C_OUTSCALAR_105_BITS(C_OUTPUT_SCALAR_105_WIDTH),
        .C_OUTSCALAR_106_BITS(C_OUTPUT_SCALAR_106_WIDTH),
        .C_OUTSCALAR_107_BITS(C_OUTPUT_SCALAR_107_WIDTH),
        .C_OUTSCALAR_108_BITS(C_OUTPUT_SCALAR_108_WIDTH),
        .C_OUTSCALAR_109_BITS(C_OUTPUT_SCALAR_109_WIDTH),
        .C_OUTSCALAR_110_BITS(C_OUTPUT_SCALAR_110_WIDTH),
        .C_OUTSCALAR_111_BITS(C_OUTPUT_SCALAR_111_WIDTH),
        .C_OUTSCALAR_112_BITS(C_OUTPUT_SCALAR_112_WIDTH),
        .C_OUTSCALAR_113_BITS(C_OUTPUT_SCALAR_113_WIDTH),
        .C_OUTSCALAR_114_BITS(C_OUTPUT_SCALAR_114_WIDTH),
        .C_OUTSCALAR_115_BITS(C_OUTPUT_SCALAR_115_WIDTH),
        .C_OUTSCALAR_116_BITS(C_OUTPUT_SCALAR_116_WIDTH),
        .C_OUTSCALAR_117_BITS(C_OUTPUT_SCALAR_117_WIDTH),
        .C_OUTSCALAR_118_BITS(C_OUTPUT_SCALAR_118_WIDTH),
        .C_OUTSCALAR_119_BITS(C_OUTPUT_SCALAR_119_WIDTH),
        .C_OUTSCALAR_120_BITS(C_OUTPUT_SCALAR_120_WIDTH),
        .C_OUTSCALAR_121_BITS(C_OUTPUT_SCALAR_121_WIDTH),
        .C_OUTSCALAR_122_BITS(C_OUTPUT_SCALAR_122_WIDTH),
        .C_OUTSCALAR_123_BITS(C_OUTPUT_SCALAR_123_WIDTH),
        .C_OUTSCALAR_124_BITS(C_OUTPUT_SCALAR_124_WIDTH),
        .C_OUTSCALAR_125_BITS(C_OUTPUT_SCALAR_125_WIDTH),
        .C_OUTSCALAR_126_BITS(C_OUTPUT_SCALAR_126_WIDTH),
        .C_OUTSCALAR_127_BITS(C_OUTPUT_SCALAR_127_WIDTH)
    ) scalar_i (
        .clk(s_axi_aclk),
        .acc_clk(aclk),
        //control interface
        .scalar_read_addr(scalar_read_addr),
        .scalar_re(scalar_re),
        .scalar_dout(scalar_dout),
        .scalar_we(scalar_we),
        .scalar_write_addr(scalar_write_addr),
        .scalar_din(scalar_din),
        .outscalar_capture(ap_done),
        .inscalar_next(inscalar_next),
        .inscalar_fifo_empty(inscalar_fifo_empty),
        .inscalar_fifo_full(inscalar_fifo_full),
        .outscalar_fifo_empty(outscalar_fifo_empty),
        .outscalar_fifo_full(outscalar_fifo_full),
        .outscalar_null_empty(outscalar_null_empty),
        .outscalar_null_dout(outscalar_null_dout),
        .outscalar_null_read(outscalar_null_read),
        //.scalar ports
        .inscalar0(ap_iscalar_0_dout),
        .inscalar1(ap_iscalar_1_dout),
        .inscalar2(ap_iscalar_2_dout),
        .inscalar3(ap_iscalar_3_dout),
        .inscalar4(ap_iscalar_4_dout),
        .inscalar5(ap_iscalar_5_dout),
        .inscalar6(ap_iscalar_6_dout),
        .inscalar7(ap_iscalar_7_dout),
        .inscalar8(ap_iscalar_8_dout),
        .inscalar9(ap_iscalar_9_dout),
        .inscalar10(ap_iscalar_10_dout),
        .inscalar11(ap_iscalar_11_dout),
        .inscalar12(ap_iscalar_12_dout),
        .inscalar13(ap_iscalar_13_dout),
        .inscalar14(ap_iscalar_14_dout),
        .inscalar15(ap_iscalar_15_dout),
        .inscalar16(ap_iscalar_16_dout),
        .inscalar17(ap_iscalar_17_dout),
        .inscalar18(ap_iscalar_18_dout),
        .inscalar19(ap_iscalar_19_dout),
        .inscalar20(ap_iscalar_20_dout),
        .inscalar21(ap_iscalar_21_dout),
        .inscalar22(ap_iscalar_22_dout),
        .inscalar23(ap_iscalar_23_dout),
        .inscalar24(ap_iscalar_24_dout),
        .inscalar25(ap_iscalar_25_dout),
        .inscalar26(ap_iscalar_26_dout),
        .inscalar27(ap_iscalar_27_dout),
        .inscalar28(ap_iscalar_28_dout),
        .inscalar29(ap_iscalar_29_dout),
        .inscalar30(ap_iscalar_30_dout),
        .inscalar31(ap_iscalar_31_dout),
        .inscalar32(ap_iscalar_32_dout),
        .inscalar33(ap_iscalar_33_dout),
        .inscalar34(ap_iscalar_34_dout),
        .inscalar35(ap_iscalar_35_dout),
        .inscalar36(ap_iscalar_36_dout),
        .inscalar37(ap_iscalar_37_dout),
        .inscalar38(ap_iscalar_38_dout),
        .inscalar39(ap_iscalar_39_dout),
        .inscalar40(ap_iscalar_40_dout),
        .inscalar41(ap_iscalar_41_dout),
        .inscalar42(ap_iscalar_42_dout),
        .inscalar43(ap_iscalar_43_dout),
        .inscalar44(ap_iscalar_44_dout),
        .inscalar45(ap_iscalar_45_dout),
        .inscalar46(ap_iscalar_46_dout),
        .inscalar47(ap_iscalar_47_dout),
        .inscalar48(ap_iscalar_48_dout),
        .inscalar49(ap_iscalar_49_dout),
        .inscalar50(ap_iscalar_50_dout),
        .inscalar51(ap_iscalar_51_dout),
        .inscalar52(ap_iscalar_52_dout),
        .inscalar53(ap_iscalar_53_dout),
        .inscalar54(ap_iscalar_54_dout),
        .inscalar55(ap_iscalar_55_dout),
        .inscalar56(ap_iscalar_56_dout),
        .inscalar57(ap_iscalar_57_dout),
        .inscalar58(ap_iscalar_58_dout),
        .inscalar59(ap_iscalar_59_dout),
        .inscalar60(ap_iscalar_60_dout),
        .inscalar61(ap_iscalar_61_dout),
        .inscalar62(ap_iscalar_62_dout),
        .inscalar63(ap_iscalar_63_dout),
        .inscalar64(ap_iscalar_64_dout),
        .inscalar65(ap_iscalar_65_dout),
        .inscalar66(ap_iscalar_66_dout),
        .inscalar67(ap_iscalar_67_dout),
        .inscalar68(ap_iscalar_68_dout),
        .inscalar69(ap_iscalar_69_dout),
        .inscalar70(ap_iscalar_70_dout),
        .inscalar71(ap_iscalar_71_dout),
        .inscalar72(ap_iscalar_72_dout),
        .inscalar73(ap_iscalar_73_dout),
        .inscalar74(ap_iscalar_74_dout),
        .inscalar75(ap_iscalar_75_dout),
        .inscalar76(ap_iscalar_76_dout),
        .inscalar77(ap_iscalar_77_dout),
        .inscalar78(ap_iscalar_78_dout),
        .inscalar79(ap_iscalar_79_dout),
        .inscalar80(ap_iscalar_80_dout),
        .inscalar81(ap_iscalar_81_dout),
        .inscalar82(ap_iscalar_82_dout),
        .inscalar83(ap_iscalar_83_dout),
        .inscalar84(ap_iscalar_84_dout),
        .inscalar85(ap_iscalar_85_dout),
        .inscalar86(ap_iscalar_86_dout),
        .inscalar87(ap_iscalar_87_dout),
        .inscalar88(ap_iscalar_88_dout),
        .inscalar89(ap_iscalar_89_dout),
        .inscalar90(ap_iscalar_90_dout),
        .inscalar91(ap_iscalar_91_dout),
        .inscalar92(ap_iscalar_92_dout),
        .inscalar93(ap_iscalar_93_dout),
        .inscalar94(ap_iscalar_94_dout),
        .inscalar95(ap_iscalar_95_dout),
        .inscalar96(ap_iscalar_96_dout),
        .inscalar97(ap_iscalar_97_dout),
        .inscalar98(ap_iscalar_98_dout),
        .inscalar99(ap_iscalar_99_dout),
        .inscalar100(ap_iscalar_100_dout),
        .inscalar101(ap_iscalar_101_dout),
        .inscalar102(ap_iscalar_102_dout),
        .inscalar103(ap_iscalar_103_dout),
        .inscalar104(ap_iscalar_104_dout),
        .inscalar105(ap_iscalar_105_dout),
        .inscalar106(ap_iscalar_106_dout),
        .inscalar107(ap_iscalar_107_dout),
        .inscalar108(ap_iscalar_108_dout),
        .inscalar109(ap_iscalar_109_dout),
        .inscalar110(ap_iscalar_110_dout),
        .inscalar111(ap_iscalar_111_dout),
        .inscalar112(ap_iscalar_112_dout),
        .inscalar113(ap_iscalar_113_dout),
        .inscalar114(ap_iscalar_114_dout),
        .inscalar115(ap_iscalar_115_dout),
        .inscalar116(ap_iscalar_116_dout),
        .inscalar117(ap_iscalar_117_dout),
        .inscalar118(ap_iscalar_118_dout),
        .inscalar119(ap_iscalar_119_dout),
        .inscalar120(ap_iscalar_120_dout),
        .inscalar121(ap_iscalar_121_dout),
        .inscalar122(ap_iscalar_122_dout),
        .inscalar123(ap_iscalar_123_dout),
        .inscalar124(ap_iscalar_124_dout),
        .inscalar125(ap_iscalar_125_dout),
        .inscalar126(ap_iscalar_126_dout),
        .inscalar127(ap_iscalar_127_dout),
        //.scalar ports
        .outscalar0(ap_oscalar_0_din),
        .outscalar1(ap_oscalar_1_din),
        .outscalar2(ap_oscalar_2_din),
        .outscalar3(ap_oscalar_3_din),
        .outscalar4(ap_oscalar_4_din),
        .outscalar5(ap_oscalar_5_din),
        .outscalar6(ap_oscalar_6_din),
        .outscalar7(ap_oscalar_7_din),
        .outscalar8(ap_oscalar_8_din),
        .outscalar9(ap_oscalar_9_din),
        .outscalar10(ap_oscalar_10_din),
        .outscalar11(ap_oscalar_11_din),
        .outscalar12(ap_oscalar_12_din),
        .outscalar13(ap_oscalar_13_din),
        .outscalar14(ap_oscalar_14_din),
        .outscalar15(ap_oscalar_15_din),
        .outscalar16(ap_oscalar_16_din),
        .outscalar17(ap_oscalar_17_din),
        .outscalar18(ap_oscalar_18_din),
        .outscalar19(ap_oscalar_19_din),
        .outscalar20(ap_oscalar_20_din),
        .outscalar21(ap_oscalar_21_din),
        .outscalar22(ap_oscalar_22_din),
        .outscalar23(ap_oscalar_23_din),
        .outscalar24(ap_oscalar_24_din),
        .outscalar25(ap_oscalar_25_din),
        .outscalar26(ap_oscalar_26_din),
        .outscalar27(ap_oscalar_27_din),
        .outscalar28(ap_oscalar_28_din),
        .outscalar29(ap_oscalar_29_din),
        .outscalar30(ap_oscalar_30_din),
        .outscalar31(ap_oscalar_31_din),
        .outscalar32(ap_oscalar_32_din),
        .outscalar33(ap_oscalar_33_din),
        .outscalar34(ap_oscalar_34_din),
        .outscalar35(ap_oscalar_35_din),
        .outscalar36(ap_oscalar_36_din),
        .outscalar37(ap_oscalar_37_din),
        .outscalar38(ap_oscalar_38_din),
        .outscalar39(ap_oscalar_39_din),
        .outscalar40(ap_oscalar_40_din),
        .outscalar41(ap_oscalar_41_din),
        .outscalar42(ap_oscalar_42_din),
        .outscalar43(ap_oscalar_43_din),
        .outscalar44(ap_oscalar_44_din),
        .outscalar45(ap_oscalar_45_din),
        .outscalar46(ap_oscalar_46_din),
        .outscalar47(ap_oscalar_47_din),
        .outscalar48(ap_oscalar_48_din),
        .outscalar49(ap_oscalar_49_din),
        .outscalar50(ap_oscalar_50_din),
        .outscalar51(ap_oscalar_51_din),
        .outscalar52(ap_oscalar_52_din),
        .outscalar53(ap_oscalar_53_din),
        .outscalar54(ap_oscalar_54_din),
        .outscalar55(ap_oscalar_55_din),
        .outscalar56(ap_oscalar_56_din),
        .outscalar57(ap_oscalar_57_din),
        .outscalar58(ap_oscalar_58_din),
        .outscalar59(ap_oscalar_59_din),
        .outscalar60(ap_oscalar_60_din),
        .outscalar61(ap_oscalar_61_din),
        .outscalar62(ap_oscalar_62_din),
        .outscalar63(ap_oscalar_63_din),
        .outscalar64(ap_oscalar_64_din),
        .outscalar65(ap_oscalar_65_din),
        .outscalar66(ap_oscalar_66_din),
        .outscalar67(ap_oscalar_67_din),
        .outscalar68(ap_oscalar_68_din),
        .outscalar69(ap_oscalar_69_din),
        .outscalar70(ap_oscalar_70_din),
        .outscalar71(ap_oscalar_71_din),
        .outscalar72(ap_oscalar_72_din),
        .outscalar73(ap_oscalar_73_din),
        .outscalar74(ap_oscalar_74_din),
        .outscalar75(ap_oscalar_75_din),
        .outscalar76(ap_oscalar_76_din),
        .outscalar77(ap_oscalar_77_din),
        .outscalar78(ap_oscalar_78_din),
        .outscalar79(ap_oscalar_79_din),
        .outscalar80(ap_oscalar_80_din),
        .outscalar81(ap_oscalar_81_din),
        .outscalar82(ap_oscalar_82_din),
        .outscalar83(ap_oscalar_83_din),
        .outscalar84(ap_oscalar_84_din),
        .outscalar85(ap_oscalar_85_din),
        .outscalar86(ap_oscalar_86_din),
        .outscalar87(ap_oscalar_87_din),
        .outscalar88(ap_oscalar_88_din),
        .outscalar89(ap_oscalar_89_din),
        .outscalar90(ap_oscalar_90_din),
        .outscalar91(ap_oscalar_91_din),
        .outscalar92(ap_oscalar_92_din),
        .outscalar93(ap_oscalar_93_din),
        .outscalar94(ap_oscalar_94_din),
        .outscalar95(ap_oscalar_95_din),
        .outscalar96(ap_oscalar_96_din),
        .outscalar97(ap_oscalar_97_din),
        .outscalar98(ap_oscalar_98_din),
        .outscalar99(ap_oscalar_99_din),
        .outscalar100(ap_oscalar_100_din),
        .outscalar101(ap_oscalar_101_din),
        .outscalar102(ap_oscalar_102_din),
        .outscalar103(ap_oscalar_103_din),
        .outscalar104(ap_oscalar_104_din),
        .outscalar105(ap_oscalar_105_din),
        .outscalar106(ap_oscalar_106_din),
        .outscalar107(ap_oscalar_107_din),
        .outscalar108(ap_oscalar_108_din),
        .outscalar109(ap_oscalar_109_din),
        .outscalar110(ap_oscalar_110_din),
        .outscalar111(ap_oscalar_111_din),
        .outscalar112(ap_oscalar_112_din),
        .outscalar113(ap_oscalar_113_din),
        .outscalar114(ap_oscalar_114_din),
        .outscalar115(ap_oscalar_115_din),
        .outscalar116(ap_oscalar_116_din),
        .outscalar117(ap_oscalar_117_din),
        .outscalar118(ap_oscalar_118_din),
        .outscalar119(ap_oscalar_119_din),
        .outscalar120(ap_oscalar_120_din),
        .outscalar121(ap_oscalar_121_din),
        .outscalar122(ap_oscalar_122_din),
        .outscalar123(ap_oscalar_123_din),
        .outscalar124(ap_oscalar_124_din),
        .outscalar125(ap_oscalar_125_din),
        .outscalar126(ap_oscalar_126_din),
        .outscalar127(ap_oscalar_127_din),
        //.scalar valid ports
        .outscalar0_vld(ap_oscalar_0_vld),
        .outscalar1_vld(ap_oscalar_1_vld),
        .outscalar2_vld(ap_oscalar_2_vld),
        .outscalar3_vld(ap_oscalar_3_vld),
        .outscalar4_vld(ap_oscalar_4_vld),
        .outscalar5_vld(ap_oscalar_5_vld),
        .outscalar6_vld(ap_oscalar_6_vld),
        .outscalar7_vld(ap_oscalar_7_vld),
        .outscalar8_vld(ap_oscalar_8_vld),
        .outscalar9_vld(ap_oscalar_9_vld),
        .outscalar10_vld(ap_oscalar_10_vld),
        .outscalar11_vld(ap_oscalar_11_vld),
        .outscalar12_vld(ap_oscalar_12_vld),
        .outscalar13_vld(ap_oscalar_13_vld),
        .outscalar14_vld(ap_oscalar_14_vld),
        .outscalar15_vld(ap_oscalar_15_vld),
        .outscalar16_vld(ap_oscalar_16_vld),
        .outscalar17_vld(ap_oscalar_17_vld),
        .outscalar18_vld(ap_oscalar_18_vld),
        .outscalar19_vld(ap_oscalar_19_vld),
        .outscalar20_vld(ap_oscalar_20_vld),
        .outscalar21_vld(ap_oscalar_21_vld),
        .outscalar22_vld(ap_oscalar_22_vld),
        .outscalar23_vld(ap_oscalar_23_vld),
        .outscalar24_vld(ap_oscalar_24_vld),
        .outscalar25_vld(ap_oscalar_25_vld),
        .outscalar26_vld(ap_oscalar_26_vld),
        .outscalar27_vld(ap_oscalar_27_vld),
        .outscalar28_vld(ap_oscalar_28_vld),
        .outscalar29_vld(ap_oscalar_29_vld),
        .outscalar30_vld(ap_oscalar_30_vld),
        .outscalar31_vld(ap_oscalar_31_vld),
        .outscalar32_vld(ap_oscalar_32_vld),
        .outscalar33_vld(ap_oscalar_33_vld),
        .outscalar34_vld(ap_oscalar_34_vld),
        .outscalar35_vld(ap_oscalar_35_vld),
        .outscalar36_vld(ap_oscalar_36_vld),
        .outscalar37_vld(ap_oscalar_37_vld),
        .outscalar38_vld(ap_oscalar_38_vld),
        .outscalar39_vld(ap_oscalar_39_vld),
        .outscalar40_vld(ap_oscalar_40_vld),
        .outscalar41_vld(ap_oscalar_41_vld),
        .outscalar42_vld(ap_oscalar_42_vld),
        .outscalar43_vld(ap_oscalar_43_vld),
        .outscalar44_vld(ap_oscalar_44_vld),
        .outscalar45_vld(ap_oscalar_45_vld),
        .outscalar46_vld(ap_oscalar_46_vld),
        .outscalar47_vld(ap_oscalar_47_vld),
        .outscalar48_vld(ap_oscalar_48_vld),
        .outscalar49_vld(ap_oscalar_49_vld),
        .outscalar50_vld(ap_oscalar_50_vld),
        .outscalar51_vld(ap_oscalar_51_vld),
        .outscalar52_vld(ap_oscalar_52_vld),
        .outscalar53_vld(ap_oscalar_53_vld),
        .outscalar54_vld(ap_oscalar_54_vld),
        .outscalar55_vld(ap_oscalar_55_vld),
        .outscalar56_vld(ap_oscalar_56_vld),
        .outscalar57_vld(ap_oscalar_57_vld),
        .outscalar58_vld(ap_oscalar_58_vld),
        .outscalar59_vld(ap_oscalar_59_vld),
        .outscalar60_vld(ap_oscalar_60_vld),
        .outscalar61_vld(ap_oscalar_61_vld),
        .outscalar62_vld(ap_oscalar_62_vld),
        .outscalar63_vld(ap_oscalar_63_vld),
        .outscalar64_vld(ap_oscalar_64_vld),
        .outscalar65_vld(ap_oscalar_65_vld),
        .outscalar66_vld(ap_oscalar_66_vld),
        .outscalar67_vld(ap_oscalar_67_vld),
        .outscalar68_vld(ap_oscalar_68_vld),
        .outscalar69_vld(ap_oscalar_69_vld),
        .outscalar70_vld(ap_oscalar_70_vld),
        .outscalar71_vld(ap_oscalar_71_vld),
        .outscalar72_vld(ap_oscalar_72_vld),
        .outscalar73_vld(ap_oscalar_73_vld),
        .outscalar74_vld(ap_oscalar_74_vld),
        .outscalar75_vld(ap_oscalar_75_vld),
        .outscalar76_vld(ap_oscalar_76_vld),
        .outscalar77_vld(ap_oscalar_77_vld),
        .outscalar78_vld(ap_oscalar_78_vld),
        .outscalar79_vld(ap_oscalar_79_vld),
        .outscalar80_vld(ap_oscalar_80_vld),
        .outscalar81_vld(ap_oscalar_81_vld),
        .outscalar82_vld(ap_oscalar_82_vld),
        .outscalar83_vld(ap_oscalar_83_vld),
        .outscalar84_vld(ap_oscalar_84_vld),
        .outscalar85_vld(ap_oscalar_85_vld),
        .outscalar86_vld(ap_oscalar_86_vld),
        .outscalar87_vld(ap_oscalar_87_vld),
        .outscalar88_vld(ap_oscalar_88_vld),
        .outscalar89_vld(ap_oscalar_89_vld),
        .outscalar90_vld(ap_oscalar_90_vld),
        .outscalar91_vld(ap_oscalar_91_vld),
        .outscalar92_vld(ap_oscalar_92_vld),
        .outscalar93_vld(ap_oscalar_93_vld),
        .outscalar94_vld(ap_oscalar_94_vld),
        .outscalar95_vld(ap_oscalar_95_vld),
        .outscalar96_vld(ap_oscalar_96_vld),
        .outscalar97_vld(ap_oscalar_97_vld),
        .outscalar98_vld(ap_oscalar_98_vld),
        .outscalar99_vld(ap_oscalar_99_vld),
        .outscalar100_vld(ap_oscalar_100_vld),
        .outscalar101_vld(ap_oscalar_101_vld),
        .outscalar102_vld(ap_oscalar_102_vld),
        .outscalar103_vld(ap_oscalar_103_vld),
        .outscalar104_vld(ap_oscalar_104_vld),
        .outscalar105_vld(ap_oscalar_105_vld),
        .outscalar106_vld(ap_oscalar_106_vld),
        .outscalar107_vld(ap_oscalar_107_vld),
        .outscalar108_vld(ap_oscalar_108_vld),
        .outscalar109_vld(ap_oscalar_109_vld),
        .outscalar110_vld(ap_oscalar_110_vld),
        .outscalar111_vld(ap_oscalar_111_vld),
        .outscalar112_vld(ap_oscalar_112_vld),
        .outscalar113_vld(ap_oscalar_113_vld),
        .outscalar114_vld(ap_oscalar_114_vld),
        .outscalar115_vld(ap_oscalar_115_vld),
        .outscalar116_vld(ap_oscalar_116_vld),
        .outscalar117_vld(ap_oscalar_117_vld),
        .outscalar118_vld(ap_oscalar_118_vld),
        .outscalar119_vld(ap_oscalar_119_vld),
        .outscalar120_vld(ap_oscalar_120_vld),
        .outscalar121_vld(ap_oscalar_121_vld),
        .outscalar122_vld(ap_oscalar_122_vld),
        .outscalar123_vld(ap_oscalar_123_vld),
        .outscalar124_vld(ap_oscalar_124_vld),
        .outscalar125_vld(ap_oscalar_125_vld),
        .outscalar126_vld(ap_oscalar_126_vld),
        .outscalar127_vld(ap_oscalar_127_vld)
    );
    
    in_fifo_args #(
        .C_NUM_INPUT_FIFOs(C_NUM_INPUT_FIFOs),
        .C_INPUT_FIFO_0_WIDTH(C_INPUT_FIFO_0_WIDTH),
        .C_INPUT_FIFO_1_WIDTH(C_INPUT_FIFO_1_WIDTH),
        .C_INPUT_FIFO_2_WIDTH(C_INPUT_FIFO_2_WIDTH),
        .C_INPUT_FIFO_3_WIDTH(C_INPUT_FIFO_3_WIDTH),
        .C_INPUT_FIFO_4_WIDTH(C_INPUT_FIFO_4_WIDTH),
        .C_INPUT_FIFO_5_WIDTH(C_INPUT_FIFO_5_WIDTH),
        .C_INPUT_FIFO_6_WIDTH(C_INPUT_FIFO_6_WIDTH),
        .C_INPUT_FIFO_7_WIDTH(C_INPUT_FIFO_7_WIDTH),
        .C_INPUT_FIFO_8_WIDTH(C_INPUT_FIFO_8_WIDTH),
        .C_INPUT_FIFO_9_WIDTH(C_INPUT_FIFO_9_WIDTH),
        .C_INPUT_FIFO_10_WIDTH(C_INPUT_FIFO_10_WIDTH),
        .C_INPUT_FIFO_11_WIDTH(C_INPUT_FIFO_11_WIDTH),
        .C_INPUT_FIFO_12_WIDTH(C_INPUT_FIFO_12_WIDTH),
        .C_INPUT_FIFO_13_WIDTH(C_INPUT_FIFO_13_WIDTH),
        .C_INPUT_FIFO_14_WIDTH(C_INPUT_FIFO_14_WIDTH),
        .C_INPUT_FIFO_15_WIDTH(C_INPUT_FIFO_15_WIDTH),
        .C_INPUT_FIFO_16_WIDTH(C_INPUT_FIFO_16_WIDTH),
        .C_INPUT_FIFO_17_WIDTH(C_INPUT_FIFO_17_WIDTH),
        .C_INPUT_FIFO_18_WIDTH(C_INPUT_FIFO_18_WIDTH),
        .C_INPUT_FIFO_19_WIDTH(C_INPUT_FIFO_19_WIDTH),
        .C_INPUT_FIFO_20_WIDTH(C_INPUT_FIFO_20_WIDTH),
        .C_INPUT_FIFO_21_WIDTH(C_INPUT_FIFO_21_WIDTH),
        .C_INPUT_FIFO_22_WIDTH(C_INPUT_FIFO_22_WIDTH),
        .C_INPUT_FIFO_23_WIDTH(C_INPUT_FIFO_23_WIDTH),
        .C_INPUT_FIFO_24_WIDTH(C_INPUT_FIFO_24_WIDTH),
        .C_INPUT_FIFO_25_WIDTH(C_INPUT_FIFO_25_WIDTH),
        .C_INPUT_FIFO_26_WIDTH(C_INPUT_FIFO_26_WIDTH),
        .C_INPUT_FIFO_27_WIDTH(C_INPUT_FIFO_27_WIDTH),
        .C_INPUT_FIFO_28_WIDTH(C_INPUT_FIFO_28_WIDTH),
        .C_INPUT_FIFO_29_WIDTH(C_INPUT_FIFO_29_WIDTH),
        .C_INPUT_FIFO_30_WIDTH(C_INPUT_FIFO_30_WIDTH),
        .C_INPUT_FIFO_31_WIDTH(C_INPUT_FIFO_31_WIDTH),
        .C_INPUT_FIFO_32_WIDTH(C_INPUT_FIFO_32_WIDTH),
        .C_INPUT_FIFO_33_WIDTH(C_INPUT_FIFO_33_WIDTH),
        .C_INPUT_FIFO_34_WIDTH(C_INPUT_FIFO_34_WIDTH),
        .C_INPUT_FIFO_35_WIDTH(C_INPUT_FIFO_35_WIDTH),
        .C_INPUT_FIFO_36_WIDTH(C_INPUT_FIFO_36_WIDTH),
        .C_INPUT_FIFO_37_WIDTH(C_INPUT_FIFO_37_WIDTH),
        .C_INPUT_FIFO_38_WIDTH(C_INPUT_FIFO_38_WIDTH),
        .C_INPUT_FIFO_39_WIDTH(C_INPUT_FIFO_39_WIDTH),
        .C_INPUT_FIFO_40_WIDTH(C_INPUT_FIFO_40_WIDTH),
        .C_INPUT_FIFO_41_WIDTH(C_INPUT_FIFO_41_WIDTH),
        .C_INPUT_FIFO_42_WIDTH(C_INPUT_FIFO_42_WIDTH),
        .C_INPUT_FIFO_43_WIDTH(C_INPUT_FIFO_43_WIDTH),
        .C_INPUT_FIFO_44_WIDTH(C_INPUT_FIFO_44_WIDTH),
        .C_INPUT_FIFO_45_WIDTH(C_INPUT_FIFO_45_WIDTH),
        .C_INPUT_FIFO_46_WIDTH(C_INPUT_FIFO_46_WIDTH),
        .C_INPUT_FIFO_47_WIDTH(C_INPUT_FIFO_47_WIDTH),
        .C_INPUT_FIFO_48_WIDTH(C_INPUT_FIFO_48_WIDTH),
        .C_INPUT_FIFO_49_WIDTH(C_INPUT_FIFO_49_WIDTH),
        .C_INPUT_FIFO_50_WIDTH(C_INPUT_FIFO_50_WIDTH),
        .C_INPUT_FIFO_51_WIDTH(C_INPUT_FIFO_51_WIDTH),
        .C_INPUT_FIFO_52_WIDTH(C_INPUT_FIFO_52_WIDTH),
        .C_INPUT_FIFO_53_WIDTH(C_INPUT_FIFO_53_WIDTH),
        .C_INPUT_FIFO_54_WIDTH(C_INPUT_FIFO_54_WIDTH),
        .C_INPUT_FIFO_55_WIDTH(C_INPUT_FIFO_55_WIDTH),
        .C_INPUT_FIFO_56_WIDTH(C_INPUT_FIFO_56_WIDTH),
        .C_INPUT_FIFO_57_WIDTH(C_INPUT_FIFO_57_WIDTH),
        .C_INPUT_FIFO_58_WIDTH(C_INPUT_FIFO_58_WIDTH),
        .C_INPUT_FIFO_59_WIDTH(C_INPUT_FIFO_59_WIDTH),
        .C_INPUT_FIFO_60_WIDTH(C_INPUT_FIFO_60_WIDTH),
        .C_INPUT_FIFO_61_WIDTH(C_INPUT_FIFO_61_WIDTH),
        .C_INPUT_FIFO_62_WIDTH(C_INPUT_FIFO_62_WIDTH),
        .C_INPUT_FIFO_63_WIDTH(C_INPUT_FIFO_63_WIDTH),
        .C_INPUT_FIFO_64_WIDTH(C_INPUT_FIFO_64_WIDTH),
        .C_INPUT_FIFO_65_WIDTH(C_INPUT_FIFO_65_WIDTH),
        .C_INPUT_FIFO_66_WIDTH(C_INPUT_FIFO_66_WIDTH),
        .C_INPUT_FIFO_67_WIDTH(C_INPUT_FIFO_67_WIDTH),
        .C_INPUT_FIFO_68_WIDTH(C_INPUT_FIFO_68_WIDTH),
        .C_INPUT_FIFO_69_WIDTH(C_INPUT_FIFO_69_WIDTH),
        .C_INPUT_FIFO_70_WIDTH(C_INPUT_FIFO_70_WIDTH),
        .C_INPUT_FIFO_71_WIDTH(C_INPUT_FIFO_71_WIDTH),
        .C_INPUT_FIFO_72_WIDTH(C_INPUT_FIFO_72_WIDTH),
        .C_INPUT_FIFO_73_WIDTH(C_INPUT_FIFO_73_WIDTH),
        .C_INPUT_FIFO_74_WIDTH(C_INPUT_FIFO_74_WIDTH),
        .C_INPUT_FIFO_75_WIDTH(C_INPUT_FIFO_75_WIDTH),
        .C_INPUT_FIFO_76_WIDTH(C_INPUT_FIFO_76_WIDTH),
        .C_INPUT_FIFO_77_WIDTH(C_INPUT_FIFO_77_WIDTH),
        .C_INPUT_FIFO_78_WIDTH(C_INPUT_FIFO_78_WIDTH),
        .C_INPUT_FIFO_79_WIDTH(C_INPUT_FIFO_79_WIDTH),
        .C_INPUT_FIFO_80_WIDTH(C_INPUT_FIFO_80_WIDTH),
        .C_INPUT_FIFO_81_WIDTH(C_INPUT_FIFO_81_WIDTH),
        .C_INPUT_FIFO_82_WIDTH(C_INPUT_FIFO_82_WIDTH),
        .C_INPUT_FIFO_83_WIDTH(C_INPUT_FIFO_83_WIDTH),
        .C_INPUT_FIFO_84_WIDTH(C_INPUT_FIFO_84_WIDTH),
        .C_INPUT_FIFO_85_WIDTH(C_INPUT_FIFO_85_WIDTH),
        .C_INPUT_FIFO_86_WIDTH(C_INPUT_FIFO_86_WIDTH),
        .C_INPUT_FIFO_87_WIDTH(C_INPUT_FIFO_87_WIDTH),
        .C_INPUT_FIFO_88_WIDTH(C_INPUT_FIFO_88_WIDTH),
        .C_INPUT_FIFO_89_WIDTH(C_INPUT_FIFO_89_WIDTH),
        .C_INPUT_FIFO_90_WIDTH(C_INPUT_FIFO_90_WIDTH),
        .C_INPUT_FIFO_91_WIDTH(C_INPUT_FIFO_91_WIDTH),
        .C_INPUT_FIFO_92_WIDTH(C_INPUT_FIFO_92_WIDTH),
        .C_INPUT_FIFO_93_WIDTH(C_INPUT_FIFO_93_WIDTH),
        .C_INPUT_FIFO_94_WIDTH(C_INPUT_FIFO_94_WIDTH),
        .C_INPUT_FIFO_95_WIDTH(C_INPUT_FIFO_95_WIDTH),
        .C_INPUT_FIFO_96_WIDTH(C_INPUT_FIFO_96_WIDTH),
        .C_INPUT_FIFO_97_WIDTH(C_INPUT_FIFO_97_WIDTH),
        .C_INPUT_FIFO_98_WIDTH(C_INPUT_FIFO_98_WIDTH),
        .C_INPUT_FIFO_99_WIDTH(C_INPUT_FIFO_99_WIDTH),
        .C_INPUT_FIFO_100_WIDTH(C_INPUT_FIFO_100_WIDTH),
        .C_INPUT_FIFO_101_WIDTH(C_INPUT_FIFO_101_WIDTH),
        .C_INPUT_FIFO_102_WIDTH(C_INPUT_FIFO_102_WIDTH),
        .C_INPUT_FIFO_103_WIDTH(C_INPUT_FIFO_103_WIDTH),
        .C_INPUT_FIFO_104_WIDTH(C_INPUT_FIFO_104_WIDTH),
        .C_INPUT_FIFO_105_WIDTH(C_INPUT_FIFO_105_WIDTH),
        .C_INPUT_FIFO_106_WIDTH(C_INPUT_FIFO_106_WIDTH),
        .C_INPUT_FIFO_107_WIDTH(C_INPUT_FIFO_107_WIDTH),
        .C_INPUT_FIFO_108_WIDTH(C_INPUT_FIFO_108_WIDTH),
        .C_INPUT_FIFO_109_WIDTH(C_INPUT_FIFO_109_WIDTH),
        .C_INPUT_FIFO_110_WIDTH(C_INPUT_FIFO_110_WIDTH),
        .C_INPUT_FIFO_111_WIDTH(C_INPUT_FIFO_111_WIDTH),
        .C_INPUT_FIFO_112_WIDTH(C_INPUT_FIFO_112_WIDTH),
        .C_INPUT_FIFO_113_WIDTH(C_INPUT_FIFO_113_WIDTH),
        .C_INPUT_FIFO_114_WIDTH(C_INPUT_FIFO_114_WIDTH),
        .C_INPUT_FIFO_115_WIDTH(C_INPUT_FIFO_115_WIDTH),
        .C_INPUT_FIFO_116_WIDTH(C_INPUT_FIFO_116_WIDTH),
        .C_INPUT_FIFO_117_WIDTH(C_INPUT_FIFO_117_WIDTH),
        .C_INPUT_FIFO_118_WIDTH(C_INPUT_FIFO_118_WIDTH),
        .C_INPUT_FIFO_119_WIDTH(C_INPUT_FIFO_119_WIDTH),
        .C_INPUT_FIFO_120_WIDTH(C_INPUT_FIFO_120_WIDTH),
        .C_INPUT_FIFO_121_WIDTH(C_INPUT_FIFO_121_WIDTH),
        .C_INPUT_FIFO_122_WIDTH(C_INPUT_FIFO_122_WIDTH),
        .C_INPUT_FIFO_123_WIDTH(C_INPUT_FIFO_123_WIDTH),
        .C_INPUT_FIFO_124_WIDTH(C_INPUT_FIFO_124_WIDTH),
        .C_INPUT_FIFO_125_WIDTH(C_INPUT_FIFO_125_WIDTH),
        .C_INPUT_FIFO_126_WIDTH(C_INPUT_FIFO_126_WIDTH),
        .C_INPUT_FIFO_127_WIDTH(C_INPUT_FIFO_127_WIDTH),
        .C_INPUT_FIFO_0_DEPTH(C_INPUT_FIFO_0_DEPTH),
        .C_INPUT_FIFO_1_DEPTH(C_INPUT_FIFO_1_DEPTH),
        .C_INPUT_FIFO_2_DEPTH(C_INPUT_FIFO_2_DEPTH),
        .C_INPUT_FIFO_3_DEPTH(C_INPUT_FIFO_3_DEPTH),
        .C_INPUT_FIFO_4_DEPTH(C_INPUT_FIFO_4_DEPTH),
        .C_INPUT_FIFO_5_DEPTH(C_INPUT_FIFO_5_DEPTH),
        .C_INPUT_FIFO_6_DEPTH(C_INPUT_FIFO_6_DEPTH),
        .C_INPUT_FIFO_7_DEPTH(C_INPUT_FIFO_7_DEPTH),
        .C_INPUT_FIFO_8_DEPTH(C_INPUT_FIFO_8_DEPTH),
        .C_INPUT_FIFO_9_DEPTH(C_INPUT_FIFO_9_DEPTH),
        .C_INPUT_FIFO_10_DEPTH(C_INPUT_FIFO_10_DEPTH),
        .C_INPUT_FIFO_11_DEPTH(C_INPUT_FIFO_11_DEPTH),
        .C_INPUT_FIFO_12_DEPTH(C_INPUT_FIFO_12_DEPTH),
        .C_INPUT_FIFO_13_DEPTH(C_INPUT_FIFO_13_DEPTH),
        .C_INPUT_FIFO_14_DEPTH(C_INPUT_FIFO_14_DEPTH),
        .C_INPUT_FIFO_15_DEPTH(C_INPUT_FIFO_15_DEPTH),
        .C_INPUT_FIFO_16_DEPTH(C_INPUT_FIFO_16_DEPTH),
        .C_INPUT_FIFO_17_DEPTH(C_INPUT_FIFO_17_DEPTH),
        .C_INPUT_FIFO_18_DEPTH(C_INPUT_FIFO_18_DEPTH),
        .C_INPUT_FIFO_19_DEPTH(C_INPUT_FIFO_19_DEPTH),
        .C_INPUT_FIFO_20_DEPTH(C_INPUT_FIFO_20_DEPTH),
        .C_INPUT_FIFO_21_DEPTH(C_INPUT_FIFO_21_DEPTH),
        .C_INPUT_FIFO_22_DEPTH(C_INPUT_FIFO_22_DEPTH),
        .C_INPUT_FIFO_23_DEPTH(C_INPUT_FIFO_23_DEPTH),
        .C_INPUT_FIFO_24_DEPTH(C_INPUT_FIFO_24_DEPTH),
        .C_INPUT_FIFO_25_DEPTH(C_INPUT_FIFO_25_DEPTH),
        .C_INPUT_FIFO_26_DEPTH(C_INPUT_FIFO_26_DEPTH),
        .C_INPUT_FIFO_27_DEPTH(C_INPUT_FIFO_27_DEPTH),
        .C_INPUT_FIFO_28_DEPTH(C_INPUT_FIFO_28_DEPTH),
        .C_INPUT_FIFO_29_DEPTH(C_INPUT_FIFO_29_DEPTH),
        .C_INPUT_FIFO_30_DEPTH(C_INPUT_FIFO_30_DEPTH),
        .C_INPUT_FIFO_31_DEPTH(C_INPUT_FIFO_31_DEPTH),
        .C_INPUT_FIFO_32_DEPTH(C_INPUT_FIFO_32_DEPTH),
        .C_INPUT_FIFO_33_DEPTH(C_INPUT_FIFO_33_DEPTH),
        .C_INPUT_FIFO_34_DEPTH(C_INPUT_FIFO_34_DEPTH),
        .C_INPUT_FIFO_35_DEPTH(C_INPUT_FIFO_35_DEPTH),
        .C_INPUT_FIFO_36_DEPTH(C_INPUT_FIFO_36_DEPTH),
        .C_INPUT_FIFO_37_DEPTH(C_INPUT_FIFO_37_DEPTH),
        .C_INPUT_FIFO_38_DEPTH(C_INPUT_FIFO_38_DEPTH),
        .C_INPUT_FIFO_39_DEPTH(C_INPUT_FIFO_39_DEPTH),
        .C_INPUT_FIFO_40_DEPTH(C_INPUT_FIFO_40_DEPTH),
        .C_INPUT_FIFO_41_DEPTH(C_INPUT_FIFO_41_DEPTH),
        .C_INPUT_FIFO_42_DEPTH(C_INPUT_FIFO_42_DEPTH),
        .C_INPUT_FIFO_43_DEPTH(C_INPUT_FIFO_43_DEPTH),
        .C_INPUT_FIFO_44_DEPTH(C_INPUT_FIFO_44_DEPTH),
        .C_INPUT_FIFO_45_DEPTH(C_INPUT_FIFO_45_DEPTH),
        .C_INPUT_FIFO_46_DEPTH(C_INPUT_FIFO_46_DEPTH),
        .C_INPUT_FIFO_47_DEPTH(C_INPUT_FIFO_47_DEPTH),
        .C_INPUT_FIFO_48_DEPTH(C_INPUT_FIFO_48_DEPTH),
        .C_INPUT_FIFO_49_DEPTH(C_INPUT_FIFO_49_DEPTH),
        .C_INPUT_FIFO_50_DEPTH(C_INPUT_FIFO_50_DEPTH),
        .C_INPUT_FIFO_51_DEPTH(C_INPUT_FIFO_51_DEPTH),
        .C_INPUT_FIFO_52_DEPTH(C_INPUT_FIFO_52_DEPTH),
        .C_INPUT_FIFO_53_DEPTH(C_INPUT_FIFO_53_DEPTH),
        .C_INPUT_FIFO_54_DEPTH(C_INPUT_FIFO_54_DEPTH),
        .C_INPUT_FIFO_55_DEPTH(C_INPUT_FIFO_55_DEPTH),
        .C_INPUT_FIFO_56_DEPTH(C_INPUT_FIFO_56_DEPTH),
        .C_INPUT_FIFO_57_DEPTH(C_INPUT_FIFO_57_DEPTH),
        .C_INPUT_FIFO_58_DEPTH(C_INPUT_FIFO_58_DEPTH),
        .C_INPUT_FIFO_59_DEPTH(C_INPUT_FIFO_59_DEPTH),
        .C_INPUT_FIFO_60_DEPTH(C_INPUT_FIFO_60_DEPTH),
        .C_INPUT_FIFO_61_DEPTH(C_INPUT_FIFO_61_DEPTH),
        .C_INPUT_FIFO_62_DEPTH(C_INPUT_FIFO_62_DEPTH),
        .C_INPUT_FIFO_63_DEPTH(C_INPUT_FIFO_63_DEPTH),
        .C_INPUT_FIFO_64_DEPTH(C_INPUT_FIFO_64_DEPTH),
        .C_INPUT_FIFO_65_DEPTH(C_INPUT_FIFO_65_DEPTH),
        .C_INPUT_FIFO_66_DEPTH(C_INPUT_FIFO_66_DEPTH),
        .C_INPUT_FIFO_67_DEPTH(C_INPUT_FIFO_67_DEPTH),
        .C_INPUT_FIFO_68_DEPTH(C_INPUT_FIFO_68_DEPTH),
        .C_INPUT_FIFO_69_DEPTH(C_INPUT_FIFO_69_DEPTH),
        .C_INPUT_FIFO_70_DEPTH(C_INPUT_FIFO_70_DEPTH),
        .C_INPUT_FIFO_71_DEPTH(C_INPUT_FIFO_71_DEPTH),
        .C_INPUT_FIFO_72_DEPTH(C_INPUT_FIFO_72_DEPTH),
        .C_INPUT_FIFO_73_DEPTH(C_INPUT_FIFO_73_DEPTH),
        .C_INPUT_FIFO_74_DEPTH(C_INPUT_FIFO_74_DEPTH),
        .C_INPUT_FIFO_75_DEPTH(C_INPUT_FIFO_75_DEPTH),
        .C_INPUT_FIFO_76_DEPTH(C_INPUT_FIFO_76_DEPTH),
        .C_INPUT_FIFO_77_DEPTH(C_INPUT_FIFO_77_DEPTH),
        .C_INPUT_FIFO_78_DEPTH(C_INPUT_FIFO_78_DEPTH),
        .C_INPUT_FIFO_79_DEPTH(C_INPUT_FIFO_79_DEPTH),
        .C_INPUT_FIFO_80_DEPTH(C_INPUT_FIFO_80_DEPTH),
        .C_INPUT_FIFO_81_DEPTH(C_INPUT_FIFO_81_DEPTH),
        .C_INPUT_FIFO_82_DEPTH(C_INPUT_FIFO_82_DEPTH),
        .C_INPUT_FIFO_83_DEPTH(C_INPUT_FIFO_83_DEPTH),
        .C_INPUT_FIFO_84_DEPTH(C_INPUT_FIFO_84_DEPTH),
        .C_INPUT_FIFO_85_DEPTH(C_INPUT_FIFO_85_DEPTH),
        .C_INPUT_FIFO_86_DEPTH(C_INPUT_FIFO_86_DEPTH),
        .C_INPUT_FIFO_87_DEPTH(C_INPUT_FIFO_87_DEPTH),
        .C_INPUT_FIFO_88_DEPTH(C_INPUT_FIFO_88_DEPTH),
        .C_INPUT_FIFO_89_DEPTH(C_INPUT_FIFO_89_DEPTH),
        .C_INPUT_FIFO_90_DEPTH(C_INPUT_FIFO_90_DEPTH),
        .C_INPUT_FIFO_91_DEPTH(C_INPUT_FIFO_91_DEPTH),
        .C_INPUT_FIFO_92_DEPTH(C_INPUT_FIFO_92_DEPTH),
        .C_INPUT_FIFO_93_DEPTH(C_INPUT_FIFO_93_DEPTH),
        .C_INPUT_FIFO_94_DEPTH(C_INPUT_FIFO_94_DEPTH),
        .C_INPUT_FIFO_95_DEPTH(C_INPUT_FIFO_95_DEPTH),
        .C_INPUT_FIFO_96_DEPTH(C_INPUT_FIFO_96_DEPTH),
        .C_INPUT_FIFO_97_DEPTH(C_INPUT_FIFO_97_DEPTH),
        .C_INPUT_FIFO_98_DEPTH(C_INPUT_FIFO_98_DEPTH),
        .C_INPUT_FIFO_99_DEPTH(C_INPUT_FIFO_99_DEPTH),
        .C_INPUT_FIFO_100_DEPTH(C_INPUT_FIFO_100_DEPTH),
        .C_INPUT_FIFO_101_DEPTH(C_INPUT_FIFO_101_DEPTH),
        .C_INPUT_FIFO_102_DEPTH(C_INPUT_FIFO_102_DEPTH),
        .C_INPUT_FIFO_103_DEPTH(C_INPUT_FIFO_103_DEPTH),
        .C_INPUT_FIFO_104_DEPTH(C_INPUT_FIFO_104_DEPTH),
        .C_INPUT_FIFO_105_DEPTH(C_INPUT_FIFO_105_DEPTH),
        .C_INPUT_FIFO_106_DEPTH(C_INPUT_FIFO_106_DEPTH),
        .C_INPUT_FIFO_107_DEPTH(C_INPUT_FIFO_107_DEPTH),
        .C_INPUT_FIFO_108_DEPTH(C_INPUT_FIFO_108_DEPTH),
        .C_INPUT_FIFO_109_DEPTH(C_INPUT_FIFO_109_DEPTH),
        .C_INPUT_FIFO_110_DEPTH(C_INPUT_FIFO_110_DEPTH),
        .C_INPUT_FIFO_111_DEPTH(C_INPUT_FIFO_111_DEPTH),
        .C_INPUT_FIFO_112_DEPTH(C_INPUT_FIFO_112_DEPTH),
        .C_INPUT_FIFO_113_DEPTH(C_INPUT_FIFO_113_DEPTH),
        .C_INPUT_FIFO_114_DEPTH(C_INPUT_FIFO_114_DEPTH),
        .C_INPUT_FIFO_115_DEPTH(C_INPUT_FIFO_115_DEPTH),
        .C_INPUT_FIFO_116_DEPTH(C_INPUT_FIFO_116_DEPTH),
        .C_INPUT_FIFO_117_DEPTH(C_INPUT_FIFO_117_DEPTH),
        .C_INPUT_FIFO_118_DEPTH(C_INPUT_FIFO_118_DEPTH),
        .C_INPUT_FIFO_119_DEPTH(C_INPUT_FIFO_119_DEPTH),
        .C_INPUT_FIFO_120_DEPTH(C_INPUT_FIFO_120_DEPTH),
        .C_INPUT_FIFO_121_DEPTH(C_INPUT_FIFO_121_DEPTH),
        .C_INPUT_FIFO_122_DEPTH(C_INPUT_FIFO_122_DEPTH),
        .C_INPUT_FIFO_123_DEPTH(C_INPUT_FIFO_123_DEPTH),
        .C_INPUT_FIFO_124_DEPTH(C_INPUT_FIFO_124_DEPTH),
        .C_INPUT_FIFO_125_DEPTH(C_INPUT_FIFO_125_DEPTH),
        .C_INPUT_FIFO_126_DEPTH(C_INPUT_FIFO_126_DEPTH),
        .C_INPUT_FIFO_127_DEPTH(C_INPUT_FIFO_127_DEPTH),
        .C_INPUT_FIFO_0_DMWIDTH(C_INPUT_FIFO_0_DMWIDTH),
        .C_INPUT_FIFO_1_DMWIDTH(C_INPUT_FIFO_1_DMWIDTH),
        .C_INPUT_FIFO_2_DMWIDTH(C_INPUT_FIFO_2_DMWIDTH),
        .C_INPUT_FIFO_3_DMWIDTH(C_INPUT_FIFO_3_DMWIDTH),
        .C_INPUT_FIFO_4_DMWIDTH(C_INPUT_FIFO_4_DMWIDTH),
        .C_INPUT_FIFO_5_DMWIDTH(C_INPUT_FIFO_5_DMWIDTH),
        .C_INPUT_FIFO_6_DMWIDTH(C_INPUT_FIFO_6_DMWIDTH),
        .C_INPUT_FIFO_7_DMWIDTH(C_INPUT_FIFO_7_DMWIDTH),
        .C_INPUT_FIFO_8_DMWIDTH(C_INPUT_FIFO_8_DMWIDTH),
        .C_INPUT_FIFO_9_DMWIDTH(C_INPUT_FIFO_9_DMWIDTH),
        .C_INPUT_FIFO_10_DMWIDTH(C_INPUT_FIFO_10_DMWIDTH),
        .C_INPUT_FIFO_11_DMWIDTH(C_INPUT_FIFO_11_DMWIDTH),
        .C_INPUT_FIFO_12_DMWIDTH(C_INPUT_FIFO_12_DMWIDTH),
        .C_INPUT_FIFO_13_DMWIDTH(C_INPUT_FIFO_13_DMWIDTH),
        .C_INPUT_FIFO_14_DMWIDTH(C_INPUT_FIFO_14_DMWIDTH),
        .C_INPUT_FIFO_15_DMWIDTH(C_INPUT_FIFO_15_DMWIDTH),
        .C_INPUT_FIFO_16_DMWIDTH(C_INPUT_FIFO_16_DMWIDTH),
        .C_INPUT_FIFO_17_DMWIDTH(C_INPUT_FIFO_17_DMWIDTH),
        .C_INPUT_FIFO_18_DMWIDTH(C_INPUT_FIFO_18_DMWIDTH),
        .C_INPUT_FIFO_19_DMWIDTH(C_INPUT_FIFO_19_DMWIDTH),
        .C_INPUT_FIFO_20_DMWIDTH(C_INPUT_FIFO_20_DMWIDTH),
        .C_INPUT_FIFO_21_DMWIDTH(C_INPUT_FIFO_21_DMWIDTH),
        .C_INPUT_FIFO_22_DMWIDTH(C_INPUT_FIFO_22_DMWIDTH),
        .C_INPUT_FIFO_23_DMWIDTH(C_INPUT_FIFO_23_DMWIDTH),
        .C_INPUT_FIFO_24_DMWIDTH(C_INPUT_FIFO_24_DMWIDTH),
        .C_INPUT_FIFO_25_DMWIDTH(C_INPUT_FIFO_25_DMWIDTH),
        .C_INPUT_FIFO_26_DMWIDTH(C_INPUT_FIFO_26_DMWIDTH),
        .C_INPUT_FIFO_27_DMWIDTH(C_INPUT_FIFO_27_DMWIDTH),
        .C_INPUT_FIFO_28_DMWIDTH(C_INPUT_FIFO_28_DMWIDTH),
        .C_INPUT_FIFO_29_DMWIDTH(C_INPUT_FIFO_29_DMWIDTH),
        .C_INPUT_FIFO_30_DMWIDTH(C_INPUT_FIFO_30_DMWIDTH),
        .C_INPUT_FIFO_31_DMWIDTH(C_INPUT_FIFO_31_DMWIDTH),
        .C_INPUT_FIFO_32_DMWIDTH(C_INPUT_FIFO_32_DMWIDTH),
        .C_INPUT_FIFO_33_DMWIDTH(C_INPUT_FIFO_33_DMWIDTH),
        .C_INPUT_FIFO_34_DMWIDTH(C_INPUT_FIFO_34_DMWIDTH),
        .C_INPUT_FIFO_35_DMWIDTH(C_INPUT_FIFO_35_DMWIDTH),
        .C_INPUT_FIFO_36_DMWIDTH(C_INPUT_FIFO_36_DMWIDTH),
        .C_INPUT_FIFO_37_DMWIDTH(C_INPUT_FIFO_37_DMWIDTH),
        .C_INPUT_FIFO_38_DMWIDTH(C_INPUT_FIFO_38_DMWIDTH),
        .C_INPUT_FIFO_39_DMWIDTH(C_INPUT_FIFO_39_DMWIDTH),
        .C_INPUT_FIFO_40_DMWIDTH(C_INPUT_FIFO_40_DMWIDTH),
        .C_INPUT_FIFO_41_DMWIDTH(C_INPUT_FIFO_41_DMWIDTH),
        .C_INPUT_FIFO_42_DMWIDTH(C_INPUT_FIFO_42_DMWIDTH),
        .C_INPUT_FIFO_43_DMWIDTH(C_INPUT_FIFO_43_DMWIDTH),
        .C_INPUT_FIFO_44_DMWIDTH(C_INPUT_FIFO_44_DMWIDTH),
        .C_INPUT_FIFO_45_DMWIDTH(C_INPUT_FIFO_45_DMWIDTH),
        .C_INPUT_FIFO_46_DMWIDTH(C_INPUT_FIFO_46_DMWIDTH),
        .C_INPUT_FIFO_47_DMWIDTH(C_INPUT_FIFO_47_DMWIDTH),
        .C_INPUT_FIFO_48_DMWIDTH(C_INPUT_FIFO_48_DMWIDTH),
        .C_INPUT_FIFO_49_DMWIDTH(C_INPUT_FIFO_49_DMWIDTH),
        .C_INPUT_FIFO_50_DMWIDTH(C_INPUT_FIFO_50_DMWIDTH),
        .C_INPUT_FIFO_51_DMWIDTH(C_INPUT_FIFO_51_DMWIDTH),
        .C_INPUT_FIFO_52_DMWIDTH(C_INPUT_FIFO_52_DMWIDTH),
        .C_INPUT_FIFO_53_DMWIDTH(C_INPUT_FIFO_53_DMWIDTH),
        .C_INPUT_FIFO_54_DMWIDTH(C_INPUT_FIFO_54_DMWIDTH),
        .C_INPUT_FIFO_55_DMWIDTH(C_INPUT_FIFO_55_DMWIDTH),
        .C_INPUT_FIFO_56_DMWIDTH(C_INPUT_FIFO_56_DMWIDTH),
        .C_INPUT_FIFO_57_DMWIDTH(C_INPUT_FIFO_57_DMWIDTH),
        .C_INPUT_FIFO_58_DMWIDTH(C_INPUT_FIFO_58_DMWIDTH),
        .C_INPUT_FIFO_59_DMWIDTH(C_INPUT_FIFO_59_DMWIDTH),
        .C_INPUT_FIFO_60_DMWIDTH(C_INPUT_FIFO_60_DMWIDTH),
        .C_INPUT_FIFO_61_DMWIDTH(C_INPUT_FIFO_61_DMWIDTH),
        .C_INPUT_FIFO_62_DMWIDTH(C_INPUT_FIFO_62_DMWIDTH),
        .C_INPUT_FIFO_63_DMWIDTH(C_INPUT_FIFO_63_DMWIDTH),
        .C_INPUT_FIFO_64_DMWIDTH(C_INPUT_FIFO_64_DMWIDTH),
        .C_INPUT_FIFO_65_DMWIDTH(C_INPUT_FIFO_65_DMWIDTH),
        .C_INPUT_FIFO_66_DMWIDTH(C_INPUT_FIFO_66_DMWIDTH),
        .C_INPUT_FIFO_67_DMWIDTH(C_INPUT_FIFO_67_DMWIDTH),
        .C_INPUT_FIFO_68_DMWIDTH(C_INPUT_FIFO_68_DMWIDTH),
        .C_INPUT_FIFO_69_DMWIDTH(C_INPUT_FIFO_69_DMWIDTH),
        .C_INPUT_FIFO_70_DMWIDTH(C_INPUT_FIFO_70_DMWIDTH),
        .C_INPUT_FIFO_71_DMWIDTH(C_INPUT_FIFO_71_DMWIDTH),
        .C_INPUT_FIFO_72_DMWIDTH(C_INPUT_FIFO_72_DMWIDTH),
        .C_INPUT_FIFO_73_DMWIDTH(C_INPUT_FIFO_73_DMWIDTH),
        .C_INPUT_FIFO_74_DMWIDTH(C_INPUT_FIFO_74_DMWIDTH),
        .C_INPUT_FIFO_75_DMWIDTH(C_INPUT_FIFO_75_DMWIDTH),
        .C_INPUT_FIFO_76_DMWIDTH(C_INPUT_FIFO_76_DMWIDTH),
        .C_INPUT_FIFO_77_DMWIDTH(C_INPUT_FIFO_77_DMWIDTH),
        .C_INPUT_FIFO_78_DMWIDTH(C_INPUT_FIFO_78_DMWIDTH),
        .C_INPUT_FIFO_79_DMWIDTH(C_INPUT_FIFO_79_DMWIDTH),
        .C_INPUT_FIFO_80_DMWIDTH(C_INPUT_FIFO_80_DMWIDTH),
        .C_INPUT_FIFO_81_DMWIDTH(C_INPUT_FIFO_81_DMWIDTH),
        .C_INPUT_FIFO_82_DMWIDTH(C_INPUT_FIFO_82_DMWIDTH),
        .C_INPUT_FIFO_83_DMWIDTH(C_INPUT_FIFO_83_DMWIDTH),
        .C_INPUT_FIFO_84_DMWIDTH(C_INPUT_FIFO_84_DMWIDTH),
        .C_INPUT_FIFO_85_DMWIDTH(C_INPUT_FIFO_85_DMWIDTH),
        .C_INPUT_FIFO_86_DMWIDTH(C_INPUT_FIFO_86_DMWIDTH),
        .C_INPUT_FIFO_87_DMWIDTH(C_INPUT_FIFO_87_DMWIDTH),
        .C_INPUT_FIFO_88_DMWIDTH(C_INPUT_FIFO_88_DMWIDTH),
        .C_INPUT_FIFO_89_DMWIDTH(C_INPUT_FIFO_89_DMWIDTH),
        .C_INPUT_FIFO_90_DMWIDTH(C_INPUT_FIFO_90_DMWIDTH),
        .C_INPUT_FIFO_91_DMWIDTH(C_INPUT_FIFO_91_DMWIDTH),
        .C_INPUT_FIFO_92_DMWIDTH(C_INPUT_FIFO_92_DMWIDTH),
        .C_INPUT_FIFO_93_DMWIDTH(C_INPUT_FIFO_93_DMWIDTH),
        .C_INPUT_FIFO_94_DMWIDTH(C_INPUT_FIFO_94_DMWIDTH),
        .C_INPUT_FIFO_95_DMWIDTH(C_INPUT_FIFO_95_DMWIDTH),
        .C_INPUT_FIFO_96_DMWIDTH(C_INPUT_FIFO_96_DMWIDTH),
        .C_INPUT_FIFO_97_DMWIDTH(C_INPUT_FIFO_97_DMWIDTH),
        .C_INPUT_FIFO_98_DMWIDTH(C_INPUT_FIFO_98_DMWIDTH),
        .C_INPUT_FIFO_99_DMWIDTH(C_INPUT_FIFO_99_DMWIDTH),
        .C_INPUT_FIFO_100_DMWIDTH(C_INPUT_FIFO_100_DMWIDTH),
        .C_INPUT_FIFO_101_DMWIDTH(C_INPUT_FIFO_101_DMWIDTH),
        .C_INPUT_FIFO_102_DMWIDTH(C_INPUT_FIFO_102_DMWIDTH),
        .C_INPUT_FIFO_103_DMWIDTH(C_INPUT_FIFO_103_DMWIDTH),
        .C_INPUT_FIFO_104_DMWIDTH(C_INPUT_FIFO_104_DMWIDTH),
        .C_INPUT_FIFO_105_DMWIDTH(C_INPUT_FIFO_105_DMWIDTH),
        .C_INPUT_FIFO_106_DMWIDTH(C_INPUT_FIFO_106_DMWIDTH),
        .C_INPUT_FIFO_107_DMWIDTH(C_INPUT_FIFO_107_DMWIDTH),
        .C_INPUT_FIFO_108_DMWIDTH(C_INPUT_FIFO_108_DMWIDTH),
        .C_INPUT_FIFO_109_DMWIDTH(C_INPUT_FIFO_109_DMWIDTH),
        .C_INPUT_FIFO_110_DMWIDTH(C_INPUT_FIFO_110_DMWIDTH),
        .C_INPUT_FIFO_111_DMWIDTH(C_INPUT_FIFO_111_DMWIDTH),
        .C_INPUT_FIFO_112_DMWIDTH(C_INPUT_FIFO_112_DMWIDTH),
        .C_INPUT_FIFO_113_DMWIDTH(C_INPUT_FIFO_113_DMWIDTH),
        .C_INPUT_FIFO_114_DMWIDTH(C_INPUT_FIFO_114_DMWIDTH),
        .C_INPUT_FIFO_115_DMWIDTH(C_INPUT_FIFO_115_DMWIDTH),
        .C_INPUT_FIFO_116_DMWIDTH(C_INPUT_FIFO_116_DMWIDTH),
        .C_INPUT_FIFO_117_DMWIDTH(C_INPUT_FIFO_117_DMWIDTH),
        .C_INPUT_FIFO_118_DMWIDTH(C_INPUT_FIFO_118_DMWIDTH),
        .C_INPUT_FIFO_119_DMWIDTH(C_INPUT_FIFO_119_DMWIDTH),
        .C_INPUT_FIFO_120_DMWIDTH(C_INPUT_FIFO_120_DMWIDTH),
        .C_INPUT_FIFO_121_DMWIDTH(C_INPUT_FIFO_121_DMWIDTH),
        .C_INPUT_FIFO_122_DMWIDTH(C_INPUT_FIFO_122_DMWIDTH),
        .C_INPUT_FIFO_123_DMWIDTH(C_INPUT_FIFO_123_DMWIDTH),
        .C_INPUT_FIFO_124_DMWIDTH(C_INPUT_FIFO_124_DMWIDTH),
        .C_INPUT_FIFO_125_DMWIDTH(C_INPUT_FIFO_125_DMWIDTH),
        .C_INPUT_FIFO_126_DMWIDTH(C_INPUT_FIFO_126_DMWIDTH),
        .C_INPUT_FIFO_127_DMWIDTH(C_INPUT_FIFO_127_DMWIDTH)
    ) in_fifo_args_i (
        .acc_clk(aclk),
        .dm_clk(s_axi_aclk),
        .aresetn(s_axi_aresetn),
        .in_fifo_allow(infifo_ctrl_allow),
        .s_axis_fifo_0_tlast(s_axis_fifo_0_tlast),
        .s_axis_fifo_0_tvalid(s_axis_fifo_0_tvalid),
        .s_axis_fifo_0_tkeep(s_axis_fifo_0_tkeep),
        .s_axis_fifo_0_tstrb(s_axis_fifo_0_tstrb),
        .s_axis_fifo_0_tdata(s_axis_fifo_0_tdata),
        .s_axis_fifo_0_tready(s_axis_fifo_0_tready),
        .ap_fifo_iarg_0_empty_n(ap_fifo_iarg_0_empty_n),
        .ap_fifo_iarg_0_dout(ap_fifo_iarg_0_dout),
        .ap_fifo_iarg_0_read(ap_fifo_iarg_0_read),
        .s_axis_fifo_1_tlast(s_axis_fifo_1_tlast),
        .s_axis_fifo_1_tvalid(s_axis_fifo_1_tvalid),
        .s_axis_fifo_1_tkeep(s_axis_fifo_1_tkeep),
        .s_axis_fifo_1_tstrb(s_axis_fifo_1_tstrb),
        .s_axis_fifo_1_tdata(s_axis_fifo_1_tdata),
        .s_axis_fifo_1_tready(s_axis_fifo_1_tready),
        .ap_fifo_iarg_1_empty_n(ap_fifo_iarg_1_empty_n),
        .ap_fifo_iarg_1_dout(ap_fifo_iarg_1_dout),
        .ap_fifo_iarg_1_read(ap_fifo_iarg_1_read),
        .s_axis_fifo_2_tlast(s_axis_fifo_2_tlast),
        .s_axis_fifo_2_tvalid(s_axis_fifo_2_tvalid),
        .s_axis_fifo_2_tkeep(s_axis_fifo_2_tkeep),
        .s_axis_fifo_2_tstrb(s_axis_fifo_2_tstrb),
        .s_axis_fifo_2_tdata(s_axis_fifo_2_tdata),
        .s_axis_fifo_2_tready(s_axis_fifo_2_tready),
        .ap_fifo_iarg_2_empty_n(ap_fifo_iarg_2_empty_n),
        .ap_fifo_iarg_2_dout(ap_fifo_iarg_2_dout),
        .ap_fifo_iarg_2_read(ap_fifo_iarg_2_read),
        .s_axis_fifo_3_tlast(s_axis_fifo_3_tlast),
        .s_axis_fifo_3_tvalid(s_axis_fifo_3_tvalid),
        .s_axis_fifo_3_tkeep(s_axis_fifo_3_tkeep),
        .s_axis_fifo_3_tstrb(s_axis_fifo_3_tstrb),
        .s_axis_fifo_3_tdata(s_axis_fifo_3_tdata),
        .s_axis_fifo_3_tready(s_axis_fifo_3_tready),
        .ap_fifo_iarg_3_empty_n(ap_fifo_iarg_3_empty_n),
        .ap_fifo_iarg_3_dout(ap_fifo_iarg_3_dout),
        .ap_fifo_iarg_3_read(ap_fifo_iarg_3_read),
        .s_axis_fifo_4_tlast(s_axis_fifo_4_tlast),
        .s_axis_fifo_4_tvalid(s_axis_fifo_4_tvalid),
        .s_axis_fifo_4_tkeep(s_axis_fifo_4_tkeep),
        .s_axis_fifo_4_tstrb(s_axis_fifo_4_tstrb),
        .s_axis_fifo_4_tdata(s_axis_fifo_4_tdata),
        .s_axis_fifo_4_tready(s_axis_fifo_4_tready),
        .ap_fifo_iarg_4_empty_n(ap_fifo_iarg_4_empty_n),
        .ap_fifo_iarg_4_dout(ap_fifo_iarg_4_dout),
        .ap_fifo_iarg_4_read(ap_fifo_iarg_4_read),
        .s_axis_fifo_5_tlast(s_axis_fifo_5_tlast),
        .s_axis_fifo_5_tvalid(s_axis_fifo_5_tvalid),
        .s_axis_fifo_5_tkeep(s_axis_fifo_5_tkeep),
        .s_axis_fifo_5_tstrb(s_axis_fifo_5_tstrb),
        .s_axis_fifo_5_tdata(s_axis_fifo_5_tdata),
        .s_axis_fifo_5_tready(s_axis_fifo_5_tready),
        .ap_fifo_iarg_5_empty_n(ap_fifo_iarg_5_empty_n),
        .ap_fifo_iarg_5_dout(ap_fifo_iarg_5_dout),
        .ap_fifo_iarg_5_read(ap_fifo_iarg_5_read),
        .s_axis_fifo_6_tlast(s_axis_fifo_6_tlast),
        .s_axis_fifo_6_tvalid(s_axis_fifo_6_tvalid),
        .s_axis_fifo_6_tkeep(s_axis_fifo_6_tkeep),
        .s_axis_fifo_6_tstrb(s_axis_fifo_6_tstrb),
        .s_axis_fifo_6_tdata(s_axis_fifo_6_tdata),
        .s_axis_fifo_6_tready(s_axis_fifo_6_tready),
        .ap_fifo_iarg_6_empty_n(ap_fifo_iarg_6_empty_n),
        .ap_fifo_iarg_6_dout(ap_fifo_iarg_6_dout),
        .ap_fifo_iarg_6_read(ap_fifo_iarg_6_read),
        .s_axis_fifo_7_tlast(s_axis_fifo_7_tlast),
        .s_axis_fifo_7_tvalid(s_axis_fifo_7_tvalid),
        .s_axis_fifo_7_tkeep(s_axis_fifo_7_tkeep),
        .s_axis_fifo_7_tstrb(s_axis_fifo_7_tstrb),
        .s_axis_fifo_7_tdata(s_axis_fifo_7_tdata),
        .s_axis_fifo_7_tready(s_axis_fifo_7_tready),
        .ap_fifo_iarg_7_empty_n(ap_fifo_iarg_7_empty_n),
        .ap_fifo_iarg_7_dout(ap_fifo_iarg_7_dout),
        .ap_fifo_iarg_7_read(ap_fifo_iarg_7_read),
        .s_axis_fifo_8_tlast(s_axis_fifo_8_tlast),
        .s_axis_fifo_8_tvalid(s_axis_fifo_8_tvalid),
        .s_axis_fifo_8_tkeep(s_axis_fifo_8_tkeep),
        .s_axis_fifo_8_tstrb(s_axis_fifo_8_tstrb),
        .s_axis_fifo_8_tdata(s_axis_fifo_8_tdata),
        .s_axis_fifo_8_tready(s_axis_fifo_8_tready),
        .ap_fifo_iarg_8_empty_n(ap_fifo_iarg_8_empty_n),
        .ap_fifo_iarg_8_dout(ap_fifo_iarg_8_dout),
        .ap_fifo_iarg_8_read(ap_fifo_iarg_8_read),
        .s_axis_fifo_9_tlast(s_axis_fifo_9_tlast),
        .s_axis_fifo_9_tvalid(s_axis_fifo_9_tvalid),
        .s_axis_fifo_9_tkeep(s_axis_fifo_9_tkeep),
        .s_axis_fifo_9_tstrb(s_axis_fifo_9_tstrb),
        .s_axis_fifo_9_tdata(s_axis_fifo_9_tdata),
        .s_axis_fifo_9_tready(s_axis_fifo_9_tready),
        .ap_fifo_iarg_9_empty_n(ap_fifo_iarg_9_empty_n),
        .ap_fifo_iarg_9_dout(ap_fifo_iarg_9_dout),
        .ap_fifo_iarg_9_read(ap_fifo_iarg_9_read),
        .s_axis_fifo_10_tlast(s_axis_fifo_10_tlast),
        .s_axis_fifo_10_tvalid(s_axis_fifo_10_tvalid),
        .s_axis_fifo_10_tkeep(s_axis_fifo_10_tkeep),
        .s_axis_fifo_10_tstrb(s_axis_fifo_10_tstrb),
        .s_axis_fifo_10_tdata(s_axis_fifo_10_tdata),
        .s_axis_fifo_10_tready(s_axis_fifo_10_tready),
        .ap_fifo_iarg_10_empty_n(ap_fifo_iarg_10_empty_n),
        .ap_fifo_iarg_10_dout(ap_fifo_iarg_10_dout),
        .ap_fifo_iarg_10_read(ap_fifo_iarg_10_read),
        .s_axis_fifo_11_tlast(s_axis_fifo_11_tlast),
        .s_axis_fifo_11_tvalid(s_axis_fifo_11_tvalid),
        .s_axis_fifo_11_tkeep(s_axis_fifo_11_tkeep),
        .s_axis_fifo_11_tstrb(s_axis_fifo_11_tstrb),
        .s_axis_fifo_11_tdata(s_axis_fifo_11_tdata),
        .s_axis_fifo_11_tready(s_axis_fifo_11_tready),
        .ap_fifo_iarg_11_empty_n(ap_fifo_iarg_11_empty_n),
        .ap_fifo_iarg_11_dout(ap_fifo_iarg_11_dout),
        .ap_fifo_iarg_11_read(ap_fifo_iarg_11_read),
        .s_axis_fifo_12_tlast(s_axis_fifo_12_tlast),
        .s_axis_fifo_12_tvalid(s_axis_fifo_12_tvalid),
        .s_axis_fifo_12_tkeep(s_axis_fifo_12_tkeep),
        .s_axis_fifo_12_tstrb(s_axis_fifo_12_tstrb),
        .s_axis_fifo_12_tdata(s_axis_fifo_12_tdata),
        .s_axis_fifo_12_tready(s_axis_fifo_12_tready),
        .ap_fifo_iarg_12_empty_n(ap_fifo_iarg_12_empty_n),
        .ap_fifo_iarg_12_dout(ap_fifo_iarg_12_dout),
        .ap_fifo_iarg_12_read(ap_fifo_iarg_12_read),
        .s_axis_fifo_13_tlast(s_axis_fifo_13_tlast),
        .s_axis_fifo_13_tvalid(s_axis_fifo_13_tvalid),
        .s_axis_fifo_13_tkeep(s_axis_fifo_13_tkeep),
        .s_axis_fifo_13_tstrb(s_axis_fifo_13_tstrb),
        .s_axis_fifo_13_tdata(s_axis_fifo_13_tdata),
        .s_axis_fifo_13_tready(s_axis_fifo_13_tready),
        .ap_fifo_iarg_13_empty_n(ap_fifo_iarg_13_empty_n),
        .ap_fifo_iarg_13_dout(ap_fifo_iarg_13_dout),
        .ap_fifo_iarg_13_read(ap_fifo_iarg_13_read),
        .s_axis_fifo_14_tlast(s_axis_fifo_14_tlast),
        .s_axis_fifo_14_tvalid(s_axis_fifo_14_tvalid),
        .s_axis_fifo_14_tkeep(s_axis_fifo_14_tkeep),
        .s_axis_fifo_14_tstrb(s_axis_fifo_14_tstrb),
        .s_axis_fifo_14_tdata(s_axis_fifo_14_tdata),
        .s_axis_fifo_14_tready(s_axis_fifo_14_tready),
        .ap_fifo_iarg_14_empty_n(ap_fifo_iarg_14_empty_n),
        .ap_fifo_iarg_14_dout(ap_fifo_iarg_14_dout),
        .ap_fifo_iarg_14_read(ap_fifo_iarg_14_read),
        .s_axis_fifo_15_tlast(s_axis_fifo_15_tlast),
        .s_axis_fifo_15_tvalid(s_axis_fifo_15_tvalid),
        .s_axis_fifo_15_tkeep(s_axis_fifo_15_tkeep),
        .s_axis_fifo_15_tstrb(s_axis_fifo_15_tstrb),
        .s_axis_fifo_15_tdata(s_axis_fifo_15_tdata),
        .s_axis_fifo_15_tready(s_axis_fifo_15_tready),
        .ap_fifo_iarg_15_empty_n(ap_fifo_iarg_15_empty_n),
        .ap_fifo_iarg_15_dout(ap_fifo_iarg_15_dout),
        .ap_fifo_iarg_15_read(ap_fifo_iarg_15_read),
        .s_axis_fifo_16_tlast(s_axis_fifo_16_tlast),
        .s_axis_fifo_16_tvalid(s_axis_fifo_16_tvalid),
        .s_axis_fifo_16_tkeep(s_axis_fifo_16_tkeep),
        .s_axis_fifo_16_tstrb(s_axis_fifo_16_tstrb),
        .s_axis_fifo_16_tdata(s_axis_fifo_16_tdata),
        .s_axis_fifo_16_tready(s_axis_fifo_16_tready),
        .ap_fifo_iarg_16_empty_n(ap_fifo_iarg_16_empty_n),
        .ap_fifo_iarg_16_dout(ap_fifo_iarg_16_dout),
        .ap_fifo_iarg_16_read(ap_fifo_iarg_16_read),
        .s_axis_fifo_17_tlast(s_axis_fifo_17_tlast),
        .s_axis_fifo_17_tvalid(s_axis_fifo_17_tvalid),
        .s_axis_fifo_17_tkeep(s_axis_fifo_17_tkeep),
        .s_axis_fifo_17_tstrb(s_axis_fifo_17_tstrb),
        .s_axis_fifo_17_tdata(s_axis_fifo_17_tdata),
        .s_axis_fifo_17_tready(s_axis_fifo_17_tready),
        .ap_fifo_iarg_17_empty_n(ap_fifo_iarg_17_empty_n),
        .ap_fifo_iarg_17_dout(ap_fifo_iarg_17_dout),
        .ap_fifo_iarg_17_read(ap_fifo_iarg_17_read),
        .s_axis_fifo_18_tlast(s_axis_fifo_18_tlast),
        .s_axis_fifo_18_tvalid(s_axis_fifo_18_tvalid),
        .s_axis_fifo_18_tkeep(s_axis_fifo_18_tkeep),
        .s_axis_fifo_18_tstrb(s_axis_fifo_18_tstrb),
        .s_axis_fifo_18_tdata(s_axis_fifo_18_tdata),
        .s_axis_fifo_18_tready(s_axis_fifo_18_tready),
        .ap_fifo_iarg_18_empty_n(ap_fifo_iarg_18_empty_n),
        .ap_fifo_iarg_18_dout(ap_fifo_iarg_18_dout),
        .ap_fifo_iarg_18_read(ap_fifo_iarg_18_read),
        .s_axis_fifo_19_tlast(s_axis_fifo_19_tlast),
        .s_axis_fifo_19_tvalid(s_axis_fifo_19_tvalid),
        .s_axis_fifo_19_tkeep(s_axis_fifo_19_tkeep),
        .s_axis_fifo_19_tstrb(s_axis_fifo_19_tstrb),
        .s_axis_fifo_19_tdata(s_axis_fifo_19_tdata),
        .s_axis_fifo_19_tready(s_axis_fifo_19_tready),
        .ap_fifo_iarg_19_empty_n(ap_fifo_iarg_19_empty_n),
        .ap_fifo_iarg_19_dout(ap_fifo_iarg_19_dout),
        .ap_fifo_iarg_19_read(ap_fifo_iarg_19_read),
        .s_axis_fifo_20_tlast(s_axis_fifo_20_tlast),
        .s_axis_fifo_20_tvalid(s_axis_fifo_20_tvalid),
        .s_axis_fifo_20_tkeep(s_axis_fifo_20_tkeep),
        .s_axis_fifo_20_tstrb(s_axis_fifo_20_tstrb),
        .s_axis_fifo_20_tdata(s_axis_fifo_20_tdata),
        .s_axis_fifo_20_tready(s_axis_fifo_20_tready),
        .ap_fifo_iarg_20_empty_n(ap_fifo_iarg_20_empty_n),
        .ap_fifo_iarg_20_dout(ap_fifo_iarg_20_dout),
        .ap_fifo_iarg_20_read(ap_fifo_iarg_20_read),
        .s_axis_fifo_21_tlast(s_axis_fifo_21_tlast),
        .s_axis_fifo_21_tvalid(s_axis_fifo_21_tvalid),
        .s_axis_fifo_21_tkeep(s_axis_fifo_21_tkeep),
        .s_axis_fifo_21_tstrb(s_axis_fifo_21_tstrb),
        .s_axis_fifo_21_tdata(s_axis_fifo_21_tdata),
        .s_axis_fifo_21_tready(s_axis_fifo_21_tready),
        .ap_fifo_iarg_21_empty_n(ap_fifo_iarg_21_empty_n),
        .ap_fifo_iarg_21_dout(ap_fifo_iarg_21_dout),
        .ap_fifo_iarg_21_read(ap_fifo_iarg_21_read),
        .s_axis_fifo_22_tlast(s_axis_fifo_22_tlast),
        .s_axis_fifo_22_tvalid(s_axis_fifo_22_tvalid),
        .s_axis_fifo_22_tkeep(s_axis_fifo_22_tkeep),
        .s_axis_fifo_22_tstrb(s_axis_fifo_22_tstrb),
        .s_axis_fifo_22_tdata(s_axis_fifo_22_tdata),
        .s_axis_fifo_22_tready(s_axis_fifo_22_tready),
        .ap_fifo_iarg_22_empty_n(ap_fifo_iarg_22_empty_n),
        .ap_fifo_iarg_22_dout(ap_fifo_iarg_22_dout),
        .ap_fifo_iarg_22_read(ap_fifo_iarg_22_read),
        .s_axis_fifo_23_tlast(s_axis_fifo_23_tlast),
        .s_axis_fifo_23_tvalid(s_axis_fifo_23_tvalid),
        .s_axis_fifo_23_tkeep(s_axis_fifo_23_tkeep),
        .s_axis_fifo_23_tstrb(s_axis_fifo_23_tstrb),
        .s_axis_fifo_23_tdata(s_axis_fifo_23_tdata),
        .s_axis_fifo_23_tready(s_axis_fifo_23_tready),
        .ap_fifo_iarg_23_empty_n(ap_fifo_iarg_23_empty_n),
        .ap_fifo_iarg_23_dout(ap_fifo_iarg_23_dout),
        .ap_fifo_iarg_23_read(ap_fifo_iarg_23_read),
        .s_axis_fifo_24_tlast(s_axis_fifo_24_tlast),
        .s_axis_fifo_24_tvalid(s_axis_fifo_24_tvalid),
        .s_axis_fifo_24_tkeep(s_axis_fifo_24_tkeep),
        .s_axis_fifo_24_tstrb(s_axis_fifo_24_tstrb),
        .s_axis_fifo_24_tdata(s_axis_fifo_24_tdata),
        .s_axis_fifo_24_tready(s_axis_fifo_24_tready),
        .ap_fifo_iarg_24_empty_n(ap_fifo_iarg_24_empty_n),
        .ap_fifo_iarg_24_dout(ap_fifo_iarg_24_dout),
        .ap_fifo_iarg_24_read(ap_fifo_iarg_24_read),
        .s_axis_fifo_25_tlast(s_axis_fifo_25_tlast),
        .s_axis_fifo_25_tvalid(s_axis_fifo_25_tvalid),
        .s_axis_fifo_25_tkeep(s_axis_fifo_25_tkeep),
        .s_axis_fifo_25_tstrb(s_axis_fifo_25_tstrb),
        .s_axis_fifo_25_tdata(s_axis_fifo_25_tdata),
        .s_axis_fifo_25_tready(s_axis_fifo_25_tready),
        .ap_fifo_iarg_25_empty_n(ap_fifo_iarg_25_empty_n),
        .ap_fifo_iarg_25_dout(ap_fifo_iarg_25_dout),
        .ap_fifo_iarg_25_read(ap_fifo_iarg_25_read),
        .s_axis_fifo_26_tlast(s_axis_fifo_26_tlast),
        .s_axis_fifo_26_tvalid(s_axis_fifo_26_tvalid),
        .s_axis_fifo_26_tkeep(s_axis_fifo_26_tkeep),
        .s_axis_fifo_26_tstrb(s_axis_fifo_26_tstrb),
        .s_axis_fifo_26_tdata(s_axis_fifo_26_tdata),
        .s_axis_fifo_26_tready(s_axis_fifo_26_tready),
        .ap_fifo_iarg_26_empty_n(ap_fifo_iarg_26_empty_n),
        .ap_fifo_iarg_26_dout(ap_fifo_iarg_26_dout),
        .ap_fifo_iarg_26_read(ap_fifo_iarg_26_read),
        .s_axis_fifo_27_tlast(s_axis_fifo_27_tlast),
        .s_axis_fifo_27_tvalid(s_axis_fifo_27_tvalid),
        .s_axis_fifo_27_tkeep(s_axis_fifo_27_tkeep),
        .s_axis_fifo_27_tstrb(s_axis_fifo_27_tstrb),
        .s_axis_fifo_27_tdata(s_axis_fifo_27_tdata),
        .s_axis_fifo_27_tready(s_axis_fifo_27_tready),
        .ap_fifo_iarg_27_empty_n(ap_fifo_iarg_27_empty_n),
        .ap_fifo_iarg_27_dout(ap_fifo_iarg_27_dout),
        .ap_fifo_iarg_27_read(ap_fifo_iarg_27_read),
        .s_axis_fifo_28_tlast(s_axis_fifo_28_tlast),
        .s_axis_fifo_28_tvalid(s_axis_fifo_28_tvalid),
        .s_axis_fifo_28_tkeep(s_axis_fifo_28_tkeep),
        .s_axis_fifo_28_tstrb(s_axis_fifo_28_tstrb),
        .s_axis_fifo_28_tdata(s_axis_fifo_28_tdata),
        .s_axis_fifo_28_tready(s_axis_fifo_28_tready),
        .ap_fifo_iarg_28_empty_n(ap_fifo_iarg_28_empty_n),
        .ap_fifo_iarg_28_dout(ap_fifo_iarg_28_dout),
        .ap_fifo_iarg_28_read(ap_fifo_iarg_28_read),
        .s_axis_fifo_29_tlast(s_axis_fifo_29_tlast),
        .s_axis_fifo_29_tvalid(s_axis_fifo_29_tvalid),
        .s_axis_fifo_29_tkeep(s_axis_fifo_29_tkeep),
        .s_axis_fifo_29_tstrb(s_axis_fifo_29_tstrb),
        .s_axis_fifo_29_tdata(s_axis_fifo_29_tdata),
        .s_axis_fifo_29_tready(s_axis_fifo_29_tready),
        .ap_fifo_iarg_29_empty_n(ap_fifo_iarg_29_empty_n),
        .ap_fifo_iarg_29_dout(ap_fifo_iarg_29_dout),
        .ap_fifo_iarg_29_read(ap_fifo_iarg_29_read),
        .s_axis_fifo_30_tlast(s_axis_fifo_30_tlast),
        .s_axis_fifo_30_tvalid(s_axis_fifo_30_tvalid),
        .s_axis_fifo_30_tkeep(s_axis_fifo_30_tkeep),
        .s_axis_fifo_30_tstrb(s_axis_fifo_30_tstrb),
        .s_axis_fifo_30_tdata(s_axis_fifo_30_tdata),
        .s_axis_fifo_30_tready(s_axis_fifo_30_tready),
        .ap_fifo_iarg_30_empty_n(ap_fifo_iarg_30_empty_n),
        .ap_fifo_iarg_30_dout(ap_fifo_iarg_30_dout),
        .ap_fifo_iarg_30_read(ap_fifo_iarg_30_read),
        .s_axis_fifo_31_tlast(s_axis_fifo_31_tlast),
        .s_axis_fifo_31_tvalid(s_axis_fifo_31_tvalid),
        .s_axis_fifo_31_tkeep(s_axis_fifo_31_tkeep),
        .s_axis_fifo_31_tstrb(s_axis_fifo_31_tstrb),
        .s_axis_fifo_31_tdata(s_axis_fifo_31_tdata),
        .s_axis_fifo_31_tready(s_axis_fifo_31_tready),
        .ap_fifo_iarg_31_empty_n(ap_fifo_iarg_31_empty_n),
        .ap_fifo_iarg_31_dout(ap_fifo_iarg_31_dout),
        .ap_fifo_iarg_31_read(ap_fifo_iarg_31_read),
        .s_axis_fifo_32_tlast(s_axis_fifo_32_tlast),
        .s_axis_fifo_32_tvalid(s_axis_fifo_32_tvalid),
        .s_axis_fifo_32_tkeep(s_axis_fifo_32_tkeep),
        .s_axis_fifo_32_tstrb(s_axis_fifo_32_tstrb),
        .s_axis_fifo_32_tdata(s_axis_fifo_32_tdata),
        .s_axis_fifo_32_tready(s_axis_fifo_32_tready),
        .ap_fifo_iarg_32_empty_n(ap_fifo_iarg_32_empty_n),
        .ap_fifo_iarg_32_dout(ap_fifo_iarg_32_dout),
        .ap_fifo_iarg_32_read(ap_fifo_iarg_32_read),
        .s_axis_fifo_33_tlast(s_axis_fifo_33_tlast),
        .s_axis_fifo_33_tvalid(s_axis_fifo_33_tvalid),
        .s_axis_fifo_33_tkeep(s_axis_fifo_33_tkeep),
        .s_axis_fifo_33_tstrb(s_axis_fifo_33_tstrb),
        .s_axis_fifo_33_tdata(s_axis_fifo_33_tdata),
        .s_axis_fifo_33_tready(s_axis_fifo_33_tready),
        .ap_fifo_iarg_33_empty_n(ap_fifo_iarg_33_empty_n),
        .ap_fifo_iarg_33_dout(ap_fifo_iarg_33_dout),
        .ap_fifo_iarg_33_read(ap_fifo_iarg_33_read),
        .s_axis_fifo_34_tlast(s_axis_fifo_34_tlast),
        .s_axis_fifo_34_tvalid(s_axis_fifo_34_tvalid),
        .s_axis_fifo_34_tkeep(s_axis_fifo_34_tkeep),
        .s_axis_fifo_34_tstrb(s_axis_fifo_34_tstrb),
        .s_axis_fifo_34_tdata(s_axis_fifo_34_tdata),
        .s_axis_fifo_34_tready(s_axis_fifo_34_tready),
        .ap_fifo_iarg_34_empty_n(ap_fifo_iarg_34_empty_n),
        .ap_fifo_iarg_34_dout(ap_fifo_iarg_34_dout),
        .ap_fifo_iarg_34_read(ap_fifo_iarg_34_read),
        .s_axis_fifo_35_tlast(s_axis_fifo_35_tlast),
        .s_axis_fifo_35_tvalid(s_axis_fifo_35_tvalid),
        .s_axis_fifo_35_tkeep(s_axis_fifo_35_tkeep),
        .s_axis_fifo_35_tstrb(s_axis_fifo_35_tstrb),
        .s_axis_fifo_35_tdata(s_axis_fifo_35_tdata),
        .s_axis_fifo_35_tready(s_axis_fifo_35_tready),
        .ap_fifo_iarg_35_empty_n(ap_fifo_iarg_35_empty_n),
        .ap_fifo_iarg_35_dout(ap_fifo_iarg_35_dout),
        .ap_fifo_iarg_35_read(ap_fifo_iarg_35_read),
        .s_axis_fifo_36_tlast(s_axis_fifo_36_tlast),
        .s_axis_fifo_36_tvalid(s_axis_fifo_36_tvalid),
        .s_axis_fifo_36_tkeep(s_axis_fifo_36_tkeep),
        .s_axis_fifo_36_tstrb(s_axis_fifo_36_tstrb),
        .s_axis_fifo_36_tdata(s_axis_fifo_36_tdata),
        .s_axis_fifo_36_tready(s_axis_fifo_36_tready),
        .ap_fifo_iarg_36_empty_n(ap_fifo_iarg_36_empty_n),
        .ap_fifo_iarg_36_dout(ap_fifo_iarg_36_dout),
        .ap_fifo_iarg_36_read(ap_fifo_iarg_36_read),
        .s_axis_fifo_37_tlast(s_axis_fifo_37_tlast),
        .s_axis_fifo_37_tvalid(s_axis_fifo_37_tvalid),
        .s_axis_fifo_37_tkeep(s_axis_fifo_37_tkeep),
        .s_axis_fifo_37_tstrb(s_axis_fifo_37_tstrb),
        .s_axis_fifo_37_tdata(s_axis_fifo_37_tdata),
        .s_axis_fifo_37_tready(s_axis_fifo_37_tready),
        .ap_fifo_iarg_37_empty_n(ap_fifo_iarg_37_empty_n),
        .ap_fifo_iarg_37_dout(ap_fifo_iarg_37_dout),
        .ap_fifo_iarg_37_read(ap_fifo_iarg_37_read),
        .s_axis_fifo_38_tlast(s_axis_fifo_38_tlast),
        .s_axis_fifo_38_tvalid(s_axis_fifo_38_tvalid),
        .s_axis_fifo_38_tkeep(s_axis_fifo_38_tkeep),
        .s_axis_fifo_38_tstrb(s_axis_fifo_38_tstrb),
        .s_axis_fifo_38_tdata(s_axis_fifo_38_tdata),
        .s_axis_fifo_38_tready(s_axis_fifo_38_tready),
        .ap_fifo_iarg_38_empty_n(ap_fifo_iarg_38_empty_n),
        .ap_fifo_iarg_38_dout(ap_fifo_iarg_38_dout),
        .ap_fifo_iarg_38_read(ap_fifo_iarg_38_read),
        .s_axis_fifo_39_tlast(s_axis_fifo_39_tlast),
        .s_axis_fifo_39_tvalid(s_axis_fifo_39_tvalid),
        .s_axis_fifo_39_tkeep(s_axis_fifo_39_tkeep),
        .s_axis_fifo_39_tstrb(s_axis_fifo_39_tstrb),
        .s_axis_fifo_39_tdata(s_axis_fifo_39_tdata),
        .s_axis_fifo_39_tready(s_axis_fifo_39_tready),
        .ap_fifo_iarg_39_empty_n(ap_fifo_iarg_39_empty_n),
        .ap_fifo_iarg_39_dout(ap_fifo_iarg_39_dout),
        .ap_fifo_iarg_39_read(ap_fifo_iarg_39_read),
        .s_axis_fifo_40_tlast(s_axis_fifo_40_tlast),
        .s_axis_fifo_40_tvalid(s_axis_fifo_40_tvalid),
        .s_axis_fifo_40_tkeep(s_axis_fifo_40_tkeep),
        .s_axis_fifo_40_tstrb(s_axis_fifo_40_tstrb),
        .s_axis_fifo_40_tdata(s_axis_fifo_40_tdata),
        .s_axis_fifo_40_tready(s_axis_fifo_40_tready),
        .ap_fifo_iarg_40_empty_n(ap_fifo_iarg_40_empty_n),
        .ap_fifo_iarg_40_dout(ap_fifo_iarg_40_dout),
        .ap_fifo_iarg_40_read(ap_fifo_iarg_40_read),
        .s_axis_fifo_41_tlast(s_axis_fifo_41_tlast),
        .s_axis_fifo_41_tvalid(s_axis_fifo_41_tvalid),
        .s_axis_fifo_41_tkeep(s_axis_fifo_41_tkeep),
        .s_axis_fifo_41_tstrb(s_axis_fifo_41_tstrb),
        .s_axis_fifo_41_tdata(s_axis_fifo_41_tdata),
        .s_axis_fifo_41_tready(s_axis_fifo_41_tready),
        .ap_fifo_iarg_41_empty_n(ap_fifo_iarg_41_empty_n),
        .ap_fifo_iarg_41_dout(ap_fifo_iarg_41_dout),
        .ap_fifo_iarg_41_read(ap_fifo_iarg_41_read),
        .s_axis_fifo_42_tlast(s_axis_fifo_42_tlast),
        .s_axis_fifo_42_tvalid(s_axis_fifo_42_tvalid),
        .s_axis_fifo_42_tkeep(s_axis_fifo_42_tkeep),
        .s_axis_fifo_42_tstrb(s_axis_fifo_42_tstrb),
        .s_axis_fifo_42_tdata(s_axis_fifo_42_tdata),
        .s_axis_fifo_42_tready(s_axis_fifo_42_tready),
        .ap_fifo_iarg_42_empty_n(ap_fifo_iarg_42_empty_n),
        .ap_fifo_iarg_42_dout(ap_fifo_iarg_42_dout),
        .ap_fifo_iarg_42_read(ap_fifo_iarg_42_read),
        .s_axis_fifo_43_tlast(s_axis_fifo_43_tlast),
        .s_axis_fifo_43_tvalid(s_axis_fifo_43_tvalid),
        .s_axis_fifo_43_tkeep(s_axis_fifo_43_tkeep),
        .s_axis_fifo_43_tstrb(s_axis_fifo_43_tstrb),
        .s_axis_fifo_43_tdata(s_axis_fifo_43_tdata),
        .s_axis_fifo_43_tready(s_axis_fifo_43_tready),
        .ap_fifo_iarg_43_empty_n(ap_fifo_iarg_43_empty_n),
        .ap_fifo_iarg_43_dout(ap_fifo_iarg_43_dout),
        .ap_fifo_iarg_43_read(ap_fifo_iarg_43_read),
        .s_axis_fifo_44_tlast(s_axis_fifo_44_tlast),
        .s_axis_fifo_44_tvalid(s_axis_fifo_44_tvalid),
        .s_axis_fifo_44_tkeep(s_axis_fifo_44_tkeep),
        .s_axis_fifo_44_tstrb(s_axis_fifo_44_tstrb),
        .s_axis_fifo_44_tdata(s_axis_fifo_44_tdata),
        .s_axis_fifo_44_tready(s_axis_fifo_44_tready),
        .ap_fifo_iarg_44_empty_n(ap_fifo_iarg_44_empty_n),
        .ap_fifo_iarg_44_dout(ap_fifo_iarg_44_dout),
        .ap_fifo_iarg_44_read(ap_fifo_iarg_44_read),
        .s_axis_fifo_45_tlast(s_axis_fifo_45_tlast),
        .s_axis_fifo_45_tvalid(s_axis_fifo_45_tvalid),
        .s_axis_fifo_45_tkeep(s_axis_fifo_45_tkeep),
        .s_axis_fifo_45_tstrb(s_axis_fifo_45_tstrb),
        .s_axis_fifo_45_tdata(s_axis_fifo_45_tdata),
        .s_axis_fifo_45_tready(s_axis_fifo_45_tready),
        .ap_fifo_iarg_45_empty_n(ap_fifo_iarg_45_empty_n),
        .ap_fifo_iarg_45_dout(ap_fifo_iarg_45_dout),
        .ap_fifo_iarg_45_read(ap_fifo_iarg_45_read),
        .s_axis_fifo_46_tlast(s_axis_fifo_46_tlast),
        .s_axis_fifo_46_tvalid(s_axis_fifo_46_tvalid),
        .s_axis_fifo_46_tkeep(s_axis_fifo_46_tkeep),
        .s_axis_fifo_46_tstrb(s_axis_fifo_46_tstrb),
        .s_axis_fifo_46_tdata(s_axis_fifo_46_tdata),
        .s_axis_fifo_46_tready(s_axis_fifo_46_tready),
        .ap_fifo_iarg_46_empty_n(ap_fifo_iarg_46_empty_n),
        .ap_fifo_iarg_46_dout(ap_fifo_iarg_46_dout),
        .ap_fifo_iarg_46_read(ap_fifo_iarg_46_read),
        .s_axis_fifo_47_tlast(s_axis_fifo_47_tlast),
        .s_axis_fifo_47_tvalid(s_axis_fifo_47_tvalid),
        .s_axis_fifo_47_tkeep(s_axis_fifo_47_tkeep),
        .s_axis_fifo_47_tstrb(s_axis_fifo_47_tstrb),
        .s_axis_fifo_47_tdata(s_axis_fifo_47_tdata),
        .s_axis_fifo_47_tready(s_axis_fifo_47_tready),
        .ap_fifo_iarg_47_empty_n(ap_fifo_iarg_47_empty_n),
        .ap_fifo_iarg_47_dout(ap_fifo_iarg_47_dout),
        .ap_fifo_iarg_47_read(ap_fifo_iarg_47_read),
        .s_axis_fifo_48_tlast(s_axis_fifo_48_tlast),
        .s_axis_fifo_48_tvalid(s_axis_fifo_48_tvalid),
        .s_axis_fifo_48_tkeep(s_axis_fifo_48_tkeep),
        .s_axis_fifo_48_tstrb(s_axis_fifo_48_tstrb),
        .s_axis_fifo_48_tdata(s_axis_fifo_48_tdata),
        .s_axis_fifo_48_tready(s_axis_fifo_48_tready),
        .ap_fifo_iarg_48_empty_n(ap_fifo_iarg_48_empty_n),
        .ap_fifo_iarg_48_dout(ap_fifo_iarg_48_dout),
        .ap_fifo_iarg_48_read(ap_fifo_iarg_48_read),
        .s_axis_fifo_49_tlast(s_axis_fifo_49_tlast),
        .s_axis_fifo_49_tvalid(s_axis_fifo_49_tvalid),
        .s_axis_fifo_49_tkeep(s_axis_fifo_49_tkeep),
        .s_axis_fifo_49_tstrb(s_axis_fifo_49_tstrb),
        .s_axis_fifo_49_tdata(s_axis_fifo_49_tdata),
        .s_axis_fifo_49_tready(s_axis_fifo_49_tready),
        .ap_fifo_iarg_49_empty_n(ap_fifo_iarg_49_empty_n),
        .ap_fifo_iarg_49_dout(ap_fifo_iarg_49_dout),
        .ap_fifo_iarg_49_read(ap_fifo_iarg_49_read),
        .s_axis_fifo_50_tlast(s_axis_fifo_50_tlast),
        .s_axis_fifo_50_tvalid(s_axis_fifo_50_tvalid),
        .s_axis_fifo_50_tkeep(s_axis_fifo_50_tkeep),
        .s_axis_fifo_50_tstrb(s_axis_fifo_50_tstrb),
        .s_axis_fifo_50_tdata(s_axis_fifo_50_tdata),
        .s_axis_fifo_50_tready(s_axis_fifo_50_tready),
        .ap_fifo_iarg_50_empty_n(ap_fifo_iarg_50_empty_n),
        .ap_fifo_iarg_50_dout(ap_fifo_iarg_50_dout),
        .ap_fifo_iarg_50_read(ap_fifo_iarg_50_read),
        .s_axis_fifo_51_tlast(s_axis_fifo_51_tlast),
        .s_axis_fifo_51_tvalid(s_axis_fifo_51_tvalid),
        .s_axis_fifo_51_tkeep(s_axis_fifo_51_tkeep),
        .s_axis_fifo_51_tstrb(s_axis_fifo_51_tstrb),
        .s_axis_fifo_51_tdata(s_axis_fifo_51_tdata),
        .s_axis_fifo_51_tready(s_axis_fifo_51_tready),
        .ap_fifo_iarg_51_empty_n(ap_fifo_iarg_51_empty_n),
        .ap_fifo_iarg_51_dout(ap_fifo_iarg_51_dout),
        .ap_fifo_iarg_51_read(ap_fifo_iarg_51_read),
        .s_axis_fifo_52_tlast(s_axis_fifo_52_tlast),
        .s_axis_fifo_52_tvalid(s_axis_fifo_52_tvalid),
        .s_axis_fifo_52_tkeep(s_axis_fifo_52_tkeep),
        .s_axis_fifo_52_tstrb(s_axis_fifo_52_tstrb),
        .s_axis_fifo_52_tdata(s_axis_fifo_52_tdata),
        .s_axis_fifo_52_tready(s_axis_fifo_52_tready),
        .ap_fifo_iarg_52_empty_n(ap_fifo_iarg_52_empty_n),
        .ap_fifo_iarg_52_dout(ap_fifo_iarg_52_dout),
        .ap_fifo_iarg_52_read(ap_fifo_iarg_52_read),
        .s_axis_fifo_53_tlast(s_axis_fifo_53_tlast),
        .s_axis_fifo_53_tvalid(s_axis_fifo_53_tvalid),
        .s_axis_fifo_53_tkeep(s_axis_fifo_53_tkeep),
        .s_axis_fifo_53_tstrb(s_axis_fifo_53_tstrb),
        .s_axis_fifo_53_tdata(s_axis_fifo_53_tdata),
        .s_axis_fifo_53_tready(s_axis_fifo_53_tready),
        .ap_fifo_iarg_53_empty_n(ap_fifo_iarg_53_empty_n),
        .ap_fifo_iarg_53_dout(ap_fifo_iarg_53_dout),
        .ap_fifo_iarg_53_read(ap_fifo_iarg_53_read),
        .s_axis_fifo_54_tlast(s_axis_fifo_54_tlast),
        .s_axis_fifo_54_tvalid(s_axis_fifo_54_tvalid),
        .s_axis_fifo_54_tkeep(s_axis_fifo_54_tkeep),
        .s_axis_fifo_54_tstrb(s_axis_fifo_54_tstrb),
        .s_axis_fifo_54_tdata(s_axis_fifo_54_tdata),
        .s_axis_fifo_54_tready(s_axis_fifo_54_tready),
        .ap_fifo_iarg_54_empty_n(ap_fifo_iarg_54_empty_n),
        .ap_fifo_iarg_54_dout(ap_fifo_iarg_54_dout),
        .ap_fifo_iarg_54_read(ap_fifo_iarg_54_read),
        .s_axis_fifo_55_tlast(s_axis_fifo_55_tlast),
        .s_axis_fifo_55_tvalid(s_axis_fifo_55_tvalid),
        .s_axis_fifo_55_tkeep(s_axis_fifo_55_tkeep),
        .s_axis_fifo_55_tstrb(s_axis_fifo_55_tstrb),
        .s_axis_fifo_55_tdata(s_axis_fifo_55_tdata),
        .s_axis_fifo_55_tready(s_axis_fifo_55_tready),
        .ap_fifo_iarg_55_empty_n(ap_fifo_iarg_55_empty_n),
        .ap_fifo_iarg_55_dout(ap_fifo_iarg_55_dout),
        .ap_fifo_iarg_55_read(ap_fifo_iarg_55_read),
        .s_axis_fifo_56_tlast(s_axis_fifo_56_tlast),
        .s_axis_fifo_56_tvalid(s_axis_fifo_56_tvalid),
        .s_axis_fifo_56_tkeep(s_axis_fifo_56_tkeep),
        .s_axis_fifo_56_tstrb(s_axis_fifo_56_tstrb),
        .s_axis_fifo_56_tdata(s_axis_fifo_56_tdata),
        .s_axis_fifo_56_tready(s_axis_fifo_56_tready),
        .ap_fifo_iarg_56_empty_n(ap_fifo_iarg_56_empty_n),
        .ap_fifo_iarg_56_dout(ap_fifo_iarg_56_dout),
        .ap_fifo_iarg_56_read(ap_fifo_iarg_56_read),
        .s_axis_fifo_57_tlast(s_axis_fifo_57_tlast),
        .s_axis_fifo_57_tvalid(s_axis_fifo_57_tvalid),
        .s_axis_fifo_57_tkeep(s_axis_fifo_57_tkeep),
        .s_axis_fifo_57_tstrb(s_axis_fifo_57_tstrb),
        .s_axis_fifo_57_tdata(s_axis_fifo_57_tdata),
        .s_axis_fifo_57_tready(s_axis_fifo_57_tready),
        .ap_fifo_iarg_57_empty_n(ap_fifo_iarg_57_empty_n),
        .ap_fifo_iarg_57_dout(ap_fifo_iarg_57_dout),
        .ap_fifo_iarg_57_read(ap_fifo_iarg_57_read),
        .s_axis_fifo_58_tlast(s_axis_fifo_58_tlast),
        .s_axis_fifo_58_tvalid(s_axis_fifo_58_tvalid),
        .s_axis_fifo_58_tkeep(s_axis_fifo_58_tkeep),
        .s_axis_fifo_58_tstrb(s_axis_fifo_58_tstrb),
        .s_axis_fifo_58_tdata(s_axis_fifo_58_tdata),
        .s_axis_fifo_58_tready(s_axis_fifo_58_tready),
        .ap_fifo_iarg_58_empty_n(ap_fifo_iarg_58_empty_n),
        .ap_fifo_iarg_58_dout(ap_fifo_iarg_58_dout),
        .ap_fifo_iarg_58_read(ap_fifo_iarg_58_read),
        .s_axis_fifo_59_tlast(s_axis_fifo_59_tlast),
        .s_axis_fifo_59_tvalid(s_axis_fifo_59_tvalid),
        .s_axis_fifo_59_tkeep(s_axis_fifo_59_tkeep),
        .s_axis_fifo_59_tstrb(s_axis_fifo_59_tstrb),
        .s_axis_fifo_59_tdata(s_axis_fifo_59_tdata),
        .s_axis_fifo_59_tready(s_axis_fifo_59_tready),
        .ap_fifo_iarg_59_empty_n(ap_fifo_iarg_59_empty_n),
        .ap_fifo_iarg_59_dout(ap_fifo_iarg_59_dout),
        .ap_fifo_iarg_59_read(ap_fifo_iarg_59_read),
        .s_axis_fifo_60_tlast(s_axis_fifo_60_tlast),
        .s_axis_fifo_60_tvalid(s_axis_fifo_60_tvalid),
        .s_axis_fifo_60_tkeep(s_axis_fifo_60_tkeep),
        .s_axis_fifo_60_tstrb(s_axis_fifo_60_tstrb),
        .s_axis_fifo_60_tdata(s_axis_fifo_60_tdata),
        .s_axis_fifo_60_tready(s_axis_fifo_60_tready),
        .ap_fifo_iarg_60_empty_n(ap_fifo_iarg_60_empty_n),
        .ap_fifo_iarg_60_dout(ap_fifo_iarg_60_dout),
        .ap_fifo_iarg_60_read(ap_fifo_iarg_60_read),
        .s_axis_fifo_61_tlast(s_axis_fifo_61_tlast),
        .s_axis_fifo_61_tvalid(s_axis_fifo_61_tvalid),
        .s_axis_fifo_61_tkeep(s_axis_fifo_61_tkeep),
        .s_axis_fifo_61_tstrb(s_axis_fifo_61_tstrb),
        .s_axis_fifo_61_tdata(s_axis_fifo_61_tdata),
        .s_axis_fifo_61_tready(s_axis_fifo_61_tready),
        .ap_fifo_iarg_61_empty_n(ap_fifo_iarg_61_empty_n),
        .ap_fifo_iarg_61_dout(ap_fifo_iarg_61_dout),
        .ap_fifo_iarg_61_read(ap_fifo_iarg_61_read),
        .s_axis_fifo_62_tlast(s_axis_fifo_62_tlast),
        .s_axis_fifo_62_tvalid(s_axis_fifo_62_tvalid),
        .s_axis_fifo_62_tkeep(s_axis_fifo_62_tkeep),
        .s_axis_fifo_62_tstrb(s_axis_fifo_62_tstrb),
        .s_axis_fifo_62_tdata(s_axis_fifo_62_tdata),
        .s_axis_fifo_62_tready(s_axis_fifo_62_tready),
        .ap_fifo_iarg_62_empty_n(ap_fifo_iarg_62_empty_n),
        .ap_fifo_iarg_62_dout(ap_fifo_iarg_62_dout),
        .ap_fifo_iarg_62_read(ap_fifo_iarg_62_read),
        .s_axis_fifo_63_tlast(s_axis_fifo_63_tlast),
        .s_axis_fifo_63_tvalid(s_axis_fifo_63_tvalid),
        .s_axis_fifo_63_tkeep(s_axis_fifo_63_tkeep),
        .s_axis_fifo_63_tstrb(s_axis_fifo_63_tstrb),
        .s_axis_fifo_63_tdata(s_axis_fifo_63_tdata),
        .s_axis_fifo_63_tready(s_axis_fifo_63_tready),
        .ap_fifo_iarg_63_empty_n(ap_fifo_iarg_63_empty_n),
        .ap_fifo_iarg_63_dout(ap_fifo_iarg_63_dout),
        .ap_fifo_iarg_63_read(ap_fifo_iarg_63_read),
        .s_axis_fifo_64_tlast(s_axis_fifo_64_tlast),
        .s_axis_fifo_64_tvalid(s_axis_fifo_64_tvalid),
        .s_axis_fifo_64_tkeep(s_axis_fifo_64_tkeep),
        .s_axis_fifo_64_tstrb(s_axis_fifo_64_tstrb),
        .s_axis_fifo_64_tdata(s_axis_fifo_64_tdata),
        .s_axis_fifo_64_tready(s_axis_fifo_64_tready),
        .ap_fifo_iarg_64_empty_n(ap_fifo_iarg_64_empty_n),
        .ap_fifo_iarg_64_dout(ap_fifo_iarg_64_dout),
        .ap_fifo_iarg_64_read(ap_fifo_iarg_64_read),
        .s_axis_fifo_65_tlast(s_axis_fifo_65_tlast),
        .s_axis_fifo_65_tvalid(s_axis_fifo_65_tvalid),
        .s_axis_fifo_65_tkeep(s_axis_fifo_65_tkeep),
        .s_axis_fifo_65_tstrb(s_axis_fifo_65_tstrb),
        .s_axis_fifo_65_tdata(s_axis_fifo_65_tdata),
        .s_axis_fifo_65_tready(s_axis_fifo_65_tready),
        .ap_fifo_iarg_65_empty_n(ap_fifo_iarg_65_empty_n),
        .ap_fifo_iarg_65_dout(ap_fifo_iarg_65_dout),
        .ap_fifo_iarg_65_read(ap_fifo_iarg_65_read),
        .s_axis_fifo_66_tlast(s_axis_fifo_66_tlast),
        .s_axis_fifo_66_tvalid(s_axis_fifo_66_tvalid),
        .s_axis_fifo_66_tkeep(s_axis_fifo_66_tkeep),
        .s_axis_fifo_66_tstrb(s_axis_fifo_66_tstrb),
        .s_axis_fifo_66_tdata(s_axis_fifo_66_tdata),
        .s_axis_fifo_66_tready(s_axis_fifo_66_tready),
        .ap_fifo_iarg_66_empty_n(ap_fifo_iarg_66_empty_n),
        .ap_fifo_iarg_66_dout(ap_fifo_iarg_66_dout),
        .ap_fifo_iarg_66_read(ap_fifo_iarg_66_read),
        .s_axis_fifo_67_tlast(s_axis_fifo_67_tlast),
        .s_axis_fifo_67_tvalid(s_axis_fifo_67_tvalid),
        .s_axis_fifo_67_tkeep(s_axis_fifo_67_tkeep),
        .s_axis_fifo_67_tstrb(s_axis_fifo_67_tstrb),
        .s_axis_fifo_67_tdata(s_axis_fifo_67_tdata),
        .s_axis_fifo_67_tready(s_axis_fifo_67_tready),
        .ap_fifo_iarg_67_empty_n(ap_fifo_iarg_67_empty_n),
        .ap_fifo_iarg_67_dout(ap_fifo_iarg_67_dout),
        .ap_fifo_iarg_67_read(ap_fifo_iarg_67_read),
        .s_axis_fifo_68_tlast(s_axis_fifo_68_tlast),
        .s_axis_fifo_68_tvalid(s_axis_fifo_68_tvalid),
        .s_axis_fifo_68_tkeep(s_axis_fifo_68_tkeep),
        .s_axis_fifo_68_tstrb(s_axis_fifo_68_tstrb),
        .s_axis_fifo_68_tdata(s_axis_fifo_68_tdata),
        .s_axis_fifo_68_tready(s_axis_fifo_68_tready),
        .ap_fifo_iarg_68_empty_n(ap_fifo_iarg_68_empty_n),
        .ap_fifo_iarg_68_dout(ap_fifo_iarg_68_dout),
        .ap_fifo_iarg_68_read(ap_fifo_iarg_68_read),
        .s_axis_fifo_69_tlast(s_axis_fifo_69_tlast),
        .s_axis_fifo_69_tvalid(s_axis_fifo_69_tvalid),
        .s_axis_fifo_69_tkeep(s_axis_fifo_69_tkeep),
        .s_axis_fifo_69_tstrb(s_axis_fifo_69_tstrb),
        .s_axis_fifo_69_tdata(s_axis_fifo_69_tdata),
        .s_axis_fifo_69_tready(s_axis_fifo_69_tready),
        .ap_fifo_iarg_69_empty_n(ap_fifo_iarg_69_empty_n),
        .ap_fifo_iarg_69_dout(ap_fifo_iarg_69_dout),
        .ap_fifo_iarg_69_read(ap_fifo_iarg_69_read),
        .s_axis_fifo_70_tlast(s_axis_fifo_70_tlast),
        .s_axis_fifo_70_tvalid(s_axis_fifo_70_tvalid),
        .s_axis_fifo_70_tkeep(s_axis_fifo_70_tkeep),
        .s_axis_fifo_70_tstrb(s_axis_fifo_70_tstrb),
        .s_axis_fifo_70_tdata(s_axis_fifo_70_tdata),
        .s_axis_fifo_70_tready(s_axis_fifo_70_tready),
        .ap_fifo_iarg_70_empty_n(ap_fifo_iarg_70_empty_n),
        .ap_fifo_iarg_70_dout(ap_fifo_iarg_70_dout),
        .ap_fifo_iarg_70_read(ap_fifo_iarg_70_read),
        .s_axis_fifo_71_tlast(s_axis_fifo_71_tlast),
        .s_axis_fifo_71_tvalid(s_axis_fifo_71_tvalid),
        .s_axis_fifo_71_tkeep(s_axis_fifo_71_tkeep),
        .s_axis_fifo_71_tstrb(s_axis_fifo_71_tstrb),
        .s_axis_fifo_71_tdata(s_axis_fifo_71_tdata),
        .s_axis_fifo_71_tready(s_axis_fifo_71_tready),
        .ap_fifo_iarg_71_empty_n(ap_fifo_iarg_71_empty_n),
        .ap_fifo_iarg_71_dout(ap_fifo_iarg_71_dout),
        .ap_fifo_iarg_71_read(ap_fifo_iarg_71_read),
        .s_axis_fifo_72_tlast(s_axis_fifo_72_tlast),
        .s_axis_fifo_72_tvalid(s_axis_fifo_72_tvalid),
        .s_axis_fifo_72_tkeep(s_axis_fifo_72_tkeep),
        .s_axis_fifo_72_tstrb(s_axis_fifo_72_tstrb),
        .s_axis_fifo_72_tdata(s_axis_fifo_72_tdata),
        .s_axis_fifo_72_tready(s_axis_fifo_72_tready),
        .ap_fifo_iarg_72_empty_n(ap_fifo_iarg_72_empty_n),
        .ap_fifo_iarg_72_dout(ap_fifo_iarg_72_dout),
        .ap_fifo_iarg_72_read(ap_fifo_iarg_72_read),
        .s_axis_fifo_73_tlast(s_axis_fifo_73_tlast),
        .s_axis_fifo_73_tvalid(s_axis_fifo_73_tvalid),
        .s_axis_fifo_73_tkeep(s_axis_fifo_73_tkeep),
        .s_axis_fifo_73_tstrb(s_axis_fifo_73_tstrb),
        .s_axis_fifo_73_tdata(s_axis_fifo_73_tdata),
        .s_axis_fifo_73_tready(s_axis_fifo_73_tready),
        .ap_fifo_iarg_73_empty_n(ap_fifo_iarg_73_empty_n),
        .ap_fifo_iarg_73_dout(ap_fifo_iarg_73_dout),
        .ap_fifo_iarg_73_read(ap_fifo_iarg_73_read),
        .s_axis_fifo_74_tlast(s_axis_fifo_74_tlast),
        .s_axis_fifo_74_tvalid(s_axis_fifo_74_tvalid),
        .s_axis_fifo_74_tkeep(s_axis_fifo_74_tkeep),
        .s_axis_fifo_74_tstrb(s_axis_fifo_74_tstrb),
        .s_axis_fifo_74_tdata(s_axis_fifo_74_tdata),
        .s_axis_fifo_74_tready(s_axis_fifo_74_tready),
        .ap_fifo_iarg_74_empty_n(ap_fifo_iarg_74_empty_n),
        .ap_fifo_iarg_74_dout(ap_fifo_iarg_74_dout),
        .ap_fifo_iarg_74_read(ap_fifo_iarg_74_read),
        .s_axis_fifo_75_tlast(s_axis_fifo_75_tlast),
        .s_axis_fifo_75_tvalid(s_axis_fifo_75_tvalid),
        .s_axis_fifo_75_tkeep(s_axis_fifo_75_tkeep),
        .s_axis_fifo_75_tstrb(s_axis_fifo_75_tstrb),
        .s_axis_fifo_75_tdata(s_axis_fifo_75_tdata),
        .s_axis_fifo_75_tready(s_axis_fifo_75_tready),
        .ap_fifo_iarg_75_empty_n(ap_fifo_iarg_75_empty_n),
        .ap_fifo_iarg_75_dout(ap_fifo_iarg_75_dout),
        .ap_fifo_iarg_75_read(ap_fifo_iarg_75_read),
        .s_axis_fifo_76_tlast(s_axis_fifo_76_tlast),
        .s_axis_fifo_76_tvalid(s_axis_fifo_76_tvalid),
        .s_axis_fifo_76_tkeep(s_axis_fifo_76_tkeep),
        .s_axis_fifo_76_tstrb(s_axis_fifo_76_tstrb),
        .s_axis_fifo_76_tdata(s_axis_fifo_76_tdata),
        .s_axis_fifo_76_tready(s_axis_fifo_76_tready),
        .ap_fifo_iarg_76_empty_n(ap_fifo_iarg_76_empty_n),
        .ap_fifo_iarg_76_dout(ap_fifo_iarg_76_dout),
        .ap_fifo_iarg_76_read(ap_fifo_iarg_76_read),
        .s_axis_fifo_77_tlast(s_axis_fifo_77_tlast),
        .s_axis_fifo_77_tvalid(s_axis_fifo_77_tvalid),
        .s_axis_fifo_77_tkeep(s_axis_fifo_77_tkeep),
        .s_axis_fifo_77_tstrb(s_axis_fifo_77_tstrb),
        .s_axis_fifo_77_tdata(s_axis_fifo_77_tdata),
        .s_axis_fifo_77_tready(s_axis_fifo_77_tready),
        .ap_fifo_iarg_77_empty_n(ap_fifo_iarg_77_empty_n),
        .ap_fifo_iarg_77_dout(ap_fifo_iarg_77_dout),
        .ap_fifo_iarg_77_read(ap_fifo_iarg_77_read),
        .s_axis_fifo_78_tlast(s_axis_fifo_78_tlast),
        .s_axis_fifo_78_tvalid(s_axis_fifo_78_tvalid),
        .s_axis_fifo_78_tkeep(s_axis_fifo_78_tkeep),
        .s_axis_fifo_78_tstrb(s_axis_fifo_78_tstrb),
        .s_axis_fifo_78_tdata(s_axis_fifo_78_tdata),
        .s_axis_fifo_78_tready(s_axis_fifo_78_tready),
        .ap_fifo_iarg_78_empty_n(ap_fifo_iarg_78_empty_n),
        .ap_fifo_iarg_78_dout(ap_fifo_iarg_78_dout),
        .ap_fifo_iarg_78_read(ap_fifo_iarg_78_read),
        .s_axis_fifo_79_tlast(s_axis_fifo_79_tlast),
        .s_axis_fifo_79_tvalid(s_axis_fifo_79_tvalid),
        .s_axis_fifo_79_tkeep(s_axis_fifo_79_tkeep),
        .s_axis_fifo_79_tstrb(s_axis_fifo_79_tstrb),
        .s_axis_fifo_79_tdata(s_axis_fifo_79_tdata),
        .s_axis_fifo_79_tready(s_axis_fifo_79_tready),
        .ap_fifo_iarg_79_empty_n(ap_fifo_iarg_79_empty_n),
        .ap_fifo_iarg_79_dout(ap_fifo_iarg_79_dout),
        .ap_fifo_iarg_79_read(ap_fifo_iarg_79_read),
        .s_axis_fifo_80_tlast(s_axis_fifo_80_tlast),
        .s_axis_fifo_80_tvalid(s_axis_fifo_80_tvalid),
        .s_axis_fifo_80_tkeep(s_axis_fifo_80_tkeep),
        .s_axis_fifo_80_tstrb(s_axis_fifo_80_tstrb),
        .s_axis_fifo_80_tdata(s_axis_fifo_80_tdata),
        .s_axis_fifo_80_tready(s_axis_fifo_80_tready),
        .ap_fifo_iarg_80_empty_n(ap_fifo_iarg_80_empty_n),
        .ap_fifo_iarg_80_dout(ap_fifo_iarg_80_dout),
        .ap_fifo_iarg_80_read(ap_fifo_iarg_80_read),
        .s_axis_fifo_81_tlast(s_axis_fifo_81_tlast),
        .s_axis_fifo_81_tvalid(s_axis_fifo_81_tvalid),
        .s_axis_fifo_81_tkeep(s_axis_fifo_81_tkeep),
        .s_axis_fifo_81_tstrb(s_axis_fifo_81_tstrb),
        .s_axis_fifo_81_tdata(s_axis_fifo_81_tdata),
        .s_axis_fifo_81_tready(s_axis_fifo_81_tready),
        .ap_fifo_iarg_81_empty_n(ap_fifo_iarg_81_empty_n),
        .ap_fifo_iarg_81_dout(ap_fifo_iarg_81_dout),
        .ap_fifo_iarg_81_read(ap_fifo_iarg_81_read),
        .s_axis_fifo_82_tlast(s_axis_fifo_82_tlast),
        .s_axis_fifo_82_tvalid(s_axis_fifo_82_tvalid),
        .s_axis_fifo_82_tkeep(s_axis_fifo_82_tkeep),
        .s_axis_fifo_82_tstrb(s_axis_fifo_82_tstrb),
        .s_axis_fifo_82_tdata(s_axis_fifo_82_tdata),
        .s_axis_fifo_82_tready(s_axis_fifo_82_tready),
        .ap_fifo_iarg_82_empty_n(ap_fifo_iarg_82_empty_n),
        .ap_fifo_iarg_82_dout(ap_fifo_iarg_82_dout),
        .ap_fifo_iarg_82_read(ap_fifo_iarg_82_read),
        .s_axis_fifo_83_tlast(s_axis_fifo_83_tlast),
        .s_axis_fifo_83_tvalid(s_axis_fifo_83_tvalid),
        .s_axis_fifo_83_tkeep(s_axis_fifo_83_tkeep),
        .s_axis_fifo_83_tstrb(s_axis_fifo_83_tstrb),
        .s_axis_fifo_83_tdata(s_axis_fifo_83_tdata),
        .s_axis_fifo_83_tready(s_axis_fifo_83_tready),
        .ap_fifo_iarg_83_empty_n(ap_fifo_iarg_83_empty_n),
        .ap_fifo_iarg_83_dout(ap_fifo_iarg_83_dout),
        .ap_fifo_iarg_83_read(ap_fifo_iarg_83_read),
        .s_axis_fifo_84_tlast(s_axis_fifo_84_tlast),
        .s_axis_fifo_84_tvalid(s_axis_fifo_84_tvalid),
        .s_axis_fifo_84_tkeep(s_axis_fifo_84_tkeep),
        .s_axis_fifo_84_tstrb(s_axis_fifo_84_tstrb),
        .s_axis_fifo_84_tdata(s_axis_fifo_84_tdata),
        .s_axis_fifo_84_tready(s_axis_fifo_84_tready),
        .ap_fifo_iarg_84_empty_n(ap_fifo_iarg_84_empty_n),
        .ap_fifo_iarg_84_dout(ap_fifo_iarg_84_dout),
        .ap_fifo_iarg_84_read(ap_fifo_iarg_84_read),
        .s_axis_fifo_85_tlast(s_axis_fifo_85_tlast),
        .s_axis_fifo_85_tvalid(s_axis_fifo_85_tvalid),
        .s_axis_fifo_85_tkeep(s_axis_fifo_85_tkeep),
        .s_axis_fifo_85_tstrb(s_axis_fifo_85_tstrb),
        .s_axis_fifo_85_tdata(s_axis_fifo_85_tdata),
        .s_axis_fifo_85_tready(s_axis_fifo_85_tready),
        .ap_fifo_iarg_85_empty_n(ap_fifo_iarg_85_empty_n),
        .ap_fifo_iarg_85_dout(ap_fifo_iarg_85_dout),
        .ap_fifo_iarg_85_read(ap_fifo_iarg_85_read),
        .s_axis_fifo_86_tlast(s_axis_fifo_86_tlast),
        .s_axis_fifo_86_tvalid(s_axis_fifo_86_tvalid),
        .s_axis_fifo_86_tkeep(s_axis_fifo_86_tkeep),
        .s_axis_fifo_86_tstrb(s_axis_fifo_86_tstrb),
        .s_axis_fifo_86_tdata(s_axis_fifo_86_tdata),
        .s_axis_fifo_86_tready(s_axis_fifo_86_tready),
        .ap_fifo_iarg_86_empty_n(ap_fifo_iarg_86_empty_n),
        .ap_fifo_iarg_86_dout(ap_fifo_iarg_86_dout),
        .ap_fifo_iarg_86_read(ap_fifo_iarg_86_read),
        .s_axis_fifo_87_tlast(s_axis_fifo_87_tlast),
        .s_axis_fifo_87_tvalid(s_axis_fifo_87_tvalid),
        .s_axis_fifo_87_tkeep(s_axis_fifo_87_tkeep),
        .s_axis_fifo_87_tstrb(s_axis_fifo_87_tstrb),
        .s_axis_fifo_87_tdata(s_axis_fifo_87_tdata),
        .s_axis_fifo_87_tready(s_axis_fifo_87_tready),
        .ap_fifo_iarg_87_empty_n(ap_fifo_iarg_87_empty_n),
        .ap_fifo_iarg_87_dout(ap_fifo_iarg_87_dout),
        .ap_fifo_iarg_87_read(ap_fifo_iarg_87_read),
        .s_axis_fifo_88_tlast(s_axis_fifo_88_tlast),
        .s_axis_fifo_88_tvalid(s_axis_fifo_88_tvalid),
        .s_axis_fifo_88_tkeep(s_axis_fifo_88_tkeep),
        .s_axis_fifo_88_tstrb(s_axis_fifo_88_tstrb),
        .s_axis_fifo_88_tdata(s_axis_fifo_88_tdata),
        .s_axis_fifo_88_tready(s_axis_fifo_88_tready),
        .ap_fifo_iarg_88_empty_n(ap_fifo_iarg_88_empty_n),
        .ap_fifo_iarg_88_dout(ap_fifo_iarg_88_dout),
        .ap_fifo_iarg_88_read(ap_fifo_iarg_88_read),
        .s_axis_fifo_89_tlast(s_axis_fifo_89_tlast),
        .s_axis_fifo_89_tvalid(s_axis_fifo_89_tvalid),
        .s_axis_fifo_89_tkeep(s_axis_fifo_89_tkeep),
        .s_axis_fifo_89_tstrb(s_axis_fifo_89_tstrb),
        .s_axis_fifo_89_tdata(s_axis_fifo_89_tdata),
        .s_axis_fifo_89_tready(s_axis_fifo_89_tready),
        .ap_fifo_iarg_89_empty_n(ap_fifo_iarg_89_empty_n),
        .ap_fifo_iarg_89_dout(ap_fifo_iarg_89_dout),
        .ap_fifo_iarg_89_read(ap_fifo_iarg_89_read),
        .s_axis_fifo_90_tlast(s_axis_fifo_90_tlast),
        .s_axis_fifo_90_tvalid(s_axis_fifo_90_tvalid),
        .s_axis_fifo_90_tkeep(s_axis_fifo_90_tkeep),
        .s_axis_fifo_90_tstrb(s_axis_fifo_90_tstrb),
        .s_axis_fifo_90_tdata(s_axis_fifo_90_tdata),
        .s_axis_fifo_90_tready(s_axis_fifo_90_tready),
        .ap_fifo_iarg_90_empty_n(ap_fifo_iarg_90_empty_n),
        .ap_fifo_iarg_90_dout(ap_fifo_iarg_90_dout),
        .ap_fifo_iarg_90_read(ap_fifo_iarg_90_read),
        .s_axis_fifo_91_tlast(s_axis_fifo_91_tlast),
        .s_axis_fifo_91_tvalid(s_axis_fifo_91_tvalid),
        .s_axis_fifo_91_tkeep(s_axis_fifo_91_tkeep),
        .s_axis_fifo_91_tstrb(s_axis_fifo_91_tstrb),
        .s_axis_fifo_91_tdata(s_axis_fifo_91_tdata),
        .s_axis_fifo_91_tready(s_axis_fifo_91_tready),
        .ap_fifo_iarg_91_empty_n(ap_fifo_iarg_91_empty_n),
        .ap_fifo_iarg_91_dout(ap_fifo_iarg_91_dout),
        .ap_fifo_iarg_91_read(ap_fifo_iarg_91_read),
        .s_axis_fifo_92_tlast(s_axis_fifo_92_tlast),
        .s_axis_fifo_92_tvalid(s_axis_fifo_92_tvalid),
        .s_axis_fifo_92_tkeep(s_axis_fifo_92_tkeep),
        .s_axis_fifo_92_tstrb(s_axis_fifo_92_tstrb),
        .s_axis_fifo_92_tdata(s_axis_fifo_92_tdata),
        .s_axis_fifo_92_tready(s_axis_fifo_92_tready),
        .ap_fifo_iarg_92_empty_n(ap_fifo_iarg_92_empty_n),
        .ap_fifo_iarg_92_dout(ap_fifo_iarg_92_dout),
        .ap_fifo_iarg_92_read(ap_fifo_iarg_92_read),
        .s_axis_fifo_93_tlast(s_axis_fifo_93_tlast),
        .s_axis_fifo_93_tvalid(s_axis_fifo_93_tvalid),
        .s_axis_fifo_93_tkeep(s_axis_fifo_93_tkeep),
        .s_axis_fifo_93_tstrb(s_axis_fifo_93_tstrb),
        .s_axis_fifo_93_tdata(s_axis_fifo_93_tdata),
        .s_axis_fifo_93_tready(s_axis_fifo_93_tready),
        .ap_fifo_iarg_93_empty_n(ap_fifo_iarg_93_empty_n),
        .ap_fifo_iarg_93_dout(ap_fifo_iarg_93_dout),
        .ap_fifo_iarg_93_read(ap_fifo_iarg_93_read),
        .s_axis_fifo_94_tlast(s_axis_fifo_94_tlast),
        .s_axis_fifo_94_tvalid(s_axis_fifo_94_tvalid),
        .s_axis_fifo_94_tkeep(s_axis_fifo_94_tkeep),
        .s_axis_fifo_94_tstrb(s_axis_fifo_94_tstrb),
        .s_axis_fifo_94_tdata(s_axis_fifo_94_tdata),
        .s_axis_fifo_94_tready(s_axis_fifo_94_tready),
        .ap_fifo_iarg_94_empty_n(ap_fifo_iarg_94_empty_n),
        .ap_fifo_iarg_94_dout(ap_fifo_iarg_94_dout),
        .ap_fifo_iarg_94_read(ap_fifo_iarg_94_read),
        .s_axis_fifo_95_tlast(s_axis_fifo_95_tlast),
        .s_axis_fifo_95_tvalid(s_axis_fifo_95_tvalid),
        .s_axis_fifo_95_tkeep(s_axis_fifo_95_tkeep),
        .s_axis_fifo_95_tstrb(s_axis_fifo_95_tstrb),
        .s_axis_fifo_95_tdata(s_axis_fifo_95_tdata),
        .s_axis_fifo_95_tready(s_axis_fifo_95_tready),
        .ap_fifo_iarg_95_empty_n(ap_fifo_iarg_95_empty_n),
        .ap_fifo_iarg_95_dout(ap_fifo_iarg_95_dout),
        .ap_fifo_iarg_95_read(ap_fifo_iarg_95_read),
        .s_axis_fifo_96_tlast(s_axis_fifo_96_tlast),
        .s_axis_fifo_96_tvalid(s_axis_fifo_96_tvalid),
        .s_axis_fifo_96_tkeep(s_axis_fifo_96_tkeep),
        .s_axis_fifo_96_tstrb(s_axis_fifo_96_tstrb),
        .s_axis_fifo_96_tdata(s_axis_fifo_96_tdata),
        .s_axis_fifo_96_tready(s_axis_fifo_96_tready),
        .ap_fifo_iarg_96_empty_n(ap_fifo_iarg_96_empty_n),
        .ap_fifo_iarg_96_dout(ap_fifo_iarg_96_dout),
        .ap_fifo_iarg_96_read(ap_fifo_iarg_96_read),
        .s_axis_fifo_97_tlast(s_axis_fifo_97_tlast),
        .s_axis_fifo_97_tvalid(s_axis_fifo_97_tvalid),
        .s_axis_fifo_97_tkeep(s_axis_fifo_97_tkeep),
        .s_axis_fifo_97_tstrb(s_axis_fifo_97_tstrb),
        .s_axis_fifo_97_tdata(s_axis_fifo_97_tdata),
        .s_axis_fifo_97_tready(s_axis_fifo_97_tready),
        .ap_fifo_iarg_97_empty_n(ap_fifo_iarg_97_empty_n),
        .ap_fifo_iarg_97_dout(ap_fifo_iarg_97_dout),
        .ap_fifo_iarg_97_read(ap_fifo_iarg_97_read),
        .s_axis_fifo_98_tlast(s_axis_fifo_98_tlast),
        .s_axis_fifo_98_tvalid(s_axis_fifo_98_tvalid),
        .s_axis_fifo_98_tkeep(s_axis_fifo_98_tkeep),
        .s_axis_fifo_98_tstrb(s_axis_fifo_98_tstrb),
        .s_axis_fifo_98_tdata(s_axis_fifo_98_tdata),
        .s_axis_fifo_98_tready(s_axis_fifo_98_tready),
        .ap_fifo_iarg_98_empty_n(ap_fifo_iarg_98_empty_n),
        .ap_fifo_iarg_98_dout(ap_fifo_iarg_98_dout),
        .ap_fifo_iarg_98_read(ap_fifo_iarg_98_read),
        .s_axis_fifo_99_tlast(s_axis_fifo_99_tlast),
        .s_axis_fifo_99_tvalid(s_axis_fifo_99_tvalid),
        .s_axis_fifo_99_tkeep(s_axis_fifo_99_tkeep),
        .s_axis_fifo_99_tstrb(s_axis_fifo_99_tstrb),
        .s_axis_fifo_99_tdata(s_axis_fifo_99_tdata),
        .s_axis_fifo_99_tready(s_axis_fifo_99_tready),
        .ap_fifo_iarg_99_empty_n(ap_fifo_iarg_99_empty_n),
        .ap_fifo_iarg_99_dout(ap_fifo_iarg_99_dout),
        .ap_fifo_iarg_99_read(ap_fifo_iarg_99_read),
        .s_axis_fifo_100_tlast(s_axis_fifo_100_tlast),
        .s_axis_fifo_100_tvalid(s_axis_fifo_100_tvalid),
        .s_axis_fifo_100_tkeep(s_axis_fifo_100_tkeep),
        .s_axis_fifo_100_tstrb(s_axis_fifo_100_tstrb),
        .s_axis_fifo_100_tdata(s_axis_fifo_100_tdata),
        .s_axis_fifo_100_tready(s_axis_fifo_100_tready),
        .ap_fifo_iarg_100_empty_n(ap_fifo_iarg_100_empty_n),
        .ap_fifo_iarg_100_dout(ap_fifo_iarg_100_dout),
        .ap_fifo_iarg_100_read(ap_fifo_iarg_100_read),
        .s_axis_fifo_101_tlast(s_axis_fifo_101_tlast),
        .s_axis_fifo_101_tvalid(s_axis_fifo_101_tvalid),
        .s_axis_fifo_101_tkeep(s_axis_fifo_101_tkeep),
        .s_axis_fifo_101_tstrb(s_axis_fifo_101_tstrb),
        .s_axis_fifo_101_tdata(s_axis_fifo_101_tdata),
        .s_axis_fifo_101_tready(s_axis_fifo_101_tready),
        .ap_fifo_iarg_101_empty_n(ap_fifo_iarg_101_empty_n),
        .ap_fifo_iarg_101_dout(ap_fifo_iarg_101_dout),
        .ap_fifo_iarg_101_read(ap_fifo_iarg_101_read),
        .s_axis_fifo_102_tlast(s_axis_fifo_102_tlast),
        .s_axis_fifo_102_tvalid(s_axis_fifo_102_tvalid),
        .s_axis_fifo_102_tkeep(s_axis_fifo_102_tkeep),
        .s_axis_fifo_102_tstrb(s_axis_fifo_102_tstrb),
        .s_axis_fifo_102_tdata(s_axis_fifo_102_tdata),
        .s_axis_fifo_102_tready(s_axis_fifo_102_tready),
        .ap_fifo_iarg_102_empty_n(ap_fifo_iarg_102_empty_n),
        .ap_fifo_iarg_102_dout(ap_fifo_iarg_102_dout),
        .ap_fifo_iarg_102_read(ap_fifo_iarg_102_read),
        .s_axis_fifo_103_tlast(s_axis_fifo_103_tlast),
        .s_axis_fifo_103_tvalid(s_axis_fifo_103_tvalid),
        .s_axis_fifo_103_tkeep(s_axis_fifo_103_tkeep),
        .s_axis_fifo_103_tstrb(s_axis_fifo_103_tstrb),
        .s_axis_fifo_103_tdata(s_axis_fifo_103_tdata),
        .s_axis_fifo_103_tready(s_axis_fifo_103_tready),
        .ap_fifo_iarg_103_empty_n(ap_fifo_iarg_103_empty_n),
        .ap_fifo_iarg_103_dout(ap_fifo_iarg_103_dout),
        .ap_fifo_iarg_103_read(ap_fifo_iarg_103_read),
        .s_axis_fifo_104_tlast(s_axis_fifo_104_tlast),
        .s_axis_fifo_104_tvalid(s_axis_fifo_104_tvalid),
        .s_axis_fifo_104_tkeep(s_axis_fifo_104_tkeep),
        .s_axis_fifo_104_tstrb(s_axis_fifo_104_tstrb),
        .s_axis_fifo_104_tdata(s_axis_fifo_104_tdata),
        .s_axis_fifo_104_tready(s_axis_fifo_104_tready),
        .ap_fifo_iarg_104_empty_n(ap_fifo_iarg_104_empty_n),
        .ap_fifo_iarg_104_dout(ap_fifo_iarg_104_dout),
        .ap_fifo_iarg_104_read(ap_fifo_iarg_104_read),
        .s_axis_fifo_105_tlast(s_axis_fifo_105_tlast),
        .s_axis_fifo_105_tvalid(s_axis_fifo_105_tvalid),
        .s_axis_fifo_105_tkeep(s_axis_fifo_105_tkeep),
        .s_axis_fifo_105_tstrb(s_axis_fifo_105_tstrb),
        .s_axis_fifo_105_tdata(s_axis_fifo_105_tdata),
        .s_axis_fifo_105_tready(s_axis_fifo_105_tready),
        .ap_fifo_iarg_105_empty_n(ap_fifo_iarg_105_empty_n),
        .ap_fifo_iarg_105_dout(ap_fifo_iarg_105_dout),
        .ap_fifo_iarg_105_read(ap_fifo_iarg_105_read),
        .s_axis_fifo_106_tlast(s_axis_fifo_106_tlast),
        .s_axis_fifo_106_tvalid(s_axis_fifo_106_tvalid),
        .s_axis_fifo_106_tkeep(s_axis_fifo_106_tkeep),
        .s_axis_fifo_106_tstrb(s_axis_fifo_106_tstrb),
        .s_axis_fifo_106_tdata(s_axis_fifo_106_tdata),
        .s_axis_fifo_106_tready(s_axis_fifo_106_tready),
        .ap_fifo_iarg_106_empty_n(ap_fifo_iarg_106_empty_n),
        .ap_fifo_iarg_106_dout(ap_fifo_iarg_106_dout),
        .ap_fifo_iarg_106_read(ap_fifo_iarg_106_read),
        .s_axis_fifo_107_tlast(s_axis_fifo_107_tlast),
        .s_axis_fifo_107_tvalid(s_axis_fifo_107_tvalid),
        .s_axis_fifo_107_tkeep(s_axis_fifo_107_tkeep),
        .s_axis_fifo_107_tstrb(s_axis_fifo_107_tstrb),
        .s_axis_fifo_107_tdata(s_axis_fifo_107_tdata),
        .s_axis_fifo_107_tready(s_axis_fifo_107_tready),
        .ap_fifo_iarg_107_empty_n(ap_fifo_iarg_107_empty_n),
        .ap_fifo_iarg_107_dout(ap_fifo_iarg_107_dout),
        .ap_fifo_iarg_107_read(ap_fifo_iarg_107_read),
        .s_axis_fifo_108_tlast(s_axis_fifo_108_tlast),
        .s_axis_fifo_108_tvalid(s_axis_fifo_108_tvalid),
        .s_axis_fifo_108_tkeep(s_axis_fifo_108_tkeep),
        .s_axis_fifo_108_tstrb(s_axis_fifo_108_tstrb),
        .s_axis_fifo_108_tdata(s_axis_fifo_108_tdata),
        .s_axis_fifo_108_tready(s_axis_fifo_108_tready),
        .ap_fifo_iarg_108_empty_n(ap_fifo_iarg_108_empty_n),
        .ap_fifo_iarg_108_dout(ap_fifo_iarg_108_dout),
        .ap_fifo_iarg_108_read(ap_fifo_iarg_108_read),
        .s_axis_fifo_109_tlast(s_axis_fifo_109_tlast),
        .s_axis_fifo_109_tvalid(s_axis_fifo_109_tvalid),
        .s_axis_fifo_109_tkeep(s_axis_fifo_109_tkeep),
        .s_axis_fifo_109_tstrb(s_axis_fifo_109_tstrb),
        .s_axis_fifo_109_tdata(s_axis_fifo_109_tdata),
        .s_axis_fifo_109_tready(s_axis_fifo_109_tready),
        .ap_fifo_iarg_109_empty_n(ap_fifo_iarg_109_empty_n),
        .ap_fifo_iarg_109_dout(ap_fifo_iarg_109_dout),
        .ap_fifo_iarg_109_read(ap_fifo_iarg_109_read),
        .s_axis_fifo_110_tlast(s_axis_fifo_110_tlast),
        .s_axis_fifo_110_tvalid(s_axis_fifo_110_tvalid),
        .s_axis_fifo_110_tkeep(s_axis_fifo_110_tkeep),
        .s_axis_fifo_110_tstrb(s_axis_fifo_110_tstrb),
        .s_axis_fifo_110_tdata(s_axis_fifo_110_tdata),
        .s_axis_fifo_110_tready(s_axis_fifo_110_tready),
        .ap_fifo_iarg_110_empty_n(ap_fifo_iarg_110_empty_n),
        .ap_fifo_iarg_110_dout(ap_fifo_iarg_110_dout),
        .ap_fifo_iarg_110_read(ap_fifo_iarg_110_read),
        .s_axis_fifo_111_tlast(s_axis_fifo_111_tlast),
        .s_axis_fifo_111_tvalid(s_axis_fifo_111_tvalid),
        .s_axis_fifo_111_tkeep(s_axis_fifo_111_tkeep),
        .s_axis_fifo_111_tstrb(s_axis_fifo_111_tstrb),
        .s_axis_fifo_111_tdata(s_axis_fifo_111_tdata),
        .s_axis_fifo_111_tready(s_axis_fifo_111_tready),
        .ap_fifo_iarg_111_empty_n(ap_fifo_iarg_111_empty_n),
        .ap_fifo_iarg_111_dout(ap_fifo_iarg_111_dout),
        .ap_fifo_iarg_111_read(ap_fifo_iarg_111_read),
        .s_axis_fifo_112_tlast(s_axis_fifo_112_tlast),
        .s_axis_fifo_112_tvalid(s_axis_fifo_112_tvalid),
        .s_axis_fifo_112_tkeep(s_axis_fifo_112_tkeep),
        .s_axis_fifo_112_tstrb(s_axis_fifo_112_tstrb),
        .s_axis_fifo_112_tdata(s_axis_fifo_112_tdata),
        .s_axis_fifo_112_tready(s_axis_fifo_112_tready),
        .ap_fifo_iarg_112_empty_n(ap_fifo_iarg_112_empty_n),
        .ap_fifo_iarg_112_dout(ap_fifo_iarg_112_dout),
        .ap_fifo_iarg_112_read(ap_fifo_iarg_112_read),
        .s_axis_fifo_113_tlast(s_axis_fifo_113_tlast),
        .s_axis_fifo_113_tvalid(s_axis_fifo_113_tvalid),
        .s_axis_fifo_113_tkeep(s_axis_fifo_113_tkeep),
        .s_axis_fifo_113_tstrb(s_axis_fifo_113_tstrb),
        .s_axis_fifo_113_tdata(s_axis_fifo_113_tdata),
        .s_axis_fifo_113_tready(s_axis_fifo_113_tready),
        .ap_fifo_iarg_113_empty_n(ap_fifo_iarg_113_empty_n),
        .ap_fifo_iarg_113_dout(ap_fifo_iarg_113_dout),
        .ap_fifo_iarg_113_read(ap_fifo_iarg_113_read),
        .s_axis_fifo_114_tlast(s_axis_fifo_114_tlast),
        .s_axis_fifo_114_tvalid(s_axis_fifo_114_tvalid),
        .s_axis_fifo_114_tkeep(s_axis_fifo_114_tkeep),
        .s_axis_fifo_114_tstrb(s_axis_fifo_114_tstrb),
        .s_axis_fifo_114_tdata(s_axis_fifo_114_tdata),
        .s_axis_fifo_114_tready(s_axis_fifo_114_tready),
        .ap_fifo_iarg_114_empty_n(ap_fifo_iarg_114_empty_n),
        .ap_fifo_iarg_114_dout(ap_fifo_iarg_114_dout),
        .ap_fifo_iarg_114_read(ap_fifo_iarg_114_read),
        .s_axis_fifo_115_tlast(s_axis_fifo_115_tlast),
        .s_axis_fifo_115_tvalid(s_axis_fifo_115_tvalid),
        .s_axis_fifo_115_tkeep(s_axis_fifo_115_tkeep),
        .s_axis_fifo_115_tstrb(s_axis_fifo_115_tstrb),
        .s_axis_fifo_115_tdata(s_axis_fifo_115_tdata),
        .s_axis_fifo_115_tready(s_axis_fifo_115_tready),
        .ap_fifo_iarg_115_empty_n(ap_fifo_iarg_115_empty_n),
        .ap_fifo_iarg_115_dout(ap_fifo_iarg_115_dout),
        .ap_fifo_iarg_115_read(ap_fifo_iarg_115_read),
        .s_axis_fifo_116_tlast(s_axis_fifo_116_tlast),
        .s_axis_fifo_116_tvalid(s_axis_fifo_116_tvalid),
        .s_axis_fifo_116_tkeep(s_axis_fifo_116_tkeep),
        .s_axis_fifo_116_tstrb(s_axis_fifo_116_tstrb),
        .s_axis_fifo_116_tdata(s_axis_fifo_116_tdata),
        .s_axis_fifo_116_tready(s_axis_fifo_116_tready),
        .ap_fifo_iarg_116_empty_n(ap_fifo_iarg_116_empty_n),
        .ap_fifo_iarg_116_dout(ap_fifo_iarg_116_dout),
        .ap_fifo_iarg_116_read(ap_fifo_iarg_116_read),
        .s_axis_fifo_117_tlast(s_axis_fifo_117_tlast),
        .s_axis_fifo_117_tvalid(s_axis_fifo_117_tvalid),
        .s_axis_fifo_117_tkeep(s_axis_fifo_117_tkeep),
        .s_axis_fifo_117_tstrb(s_axis_fifo_117_tstrb),
        .s_axis_fifo_117_tdata(s_axis_fifo_117_tdata),
        .s_axis_fifo_117_tready(s_axis_fifo_117_tready),
        .ap_fifo_iarg_117_empty_n(ap_fifo_iarg_117_empty_n),
        .ap_fifo_iarg_117_dout(ap_fifo_iarg_117_dout),
        .ap_fifo_iarg_117_read(ap_fifo_iarg_117_read),
        .s_axis_fifo_118_tlast(s_axis_fifo_118_tlast),
        .s_axis_fifo_118_tvalid(s_axis_fifo_118_tvalid),
        .s_axis_fifo_118_tkeep(s_axis_fifo_118_tkeep),
        .s_axis_fifo_118_tstrb(s_axis_fifo_118_tstrb),
        .s_axis_fifo_118_tdata(s_axis_fifo_118_tdata),
        .s_axis_fifo_118_tready(s_axis_fifo_118_tready),
        .ap_fifo_iarg_118_empty_n(ap_fifo_iarg_118_empty_n),
        .ap_fifo_iarg_118_dout(ap_fifo_iarg_118_dout),
        .ap_fifo_iarg_118_read(ap_fifo_iarg_118_read),
        .s_axis_fifo_119_tlast(s_axis_fifo_119_tlast),
        .s_axis_fifo_119_tvalid(s_axis_fifo_119_tvalid),
        .s_axis_fifo_119_tkeep(s_axis_fifo_119_tkeep),
        .s_axis_fifo_119_tstrb(s_axis_fifo_119_tstrb),
        .s_axis_fifo_119_tdata(s_axis_fifo_119_tdata),
        .s_axis_fifo_119_tready(s_axis_fifo_119_tready),
        .ap_fifo_iarg_119_empty_n(ap_fifo_iarg_119_empty_n),
        .ap_fifo_iarg_119_dout(ap_fifo_iarg_119_dout),
        .ap_fifo_iarg_119_read(ap_fifo_iarg_119_read),
        .s_axis_fifo_120_tlast(s_axis_fifo_120_tlast),
        .s_axis_fifo_120_tvalid(s_axis_fifo_120_tvalid),
        .s_axis_fifo_120_tkeep(s_axis_fifo_120_tkeep),
        .s_axis_fifo_120_tstrb(s_axis_fifo_120_tstrb),
        .s_axis_fifo_120_tdata(s_axis_fifo_120_tdata),
        .s_axis_fifo_120_tready(s_axis_fifo_120_tready),
        .ap_fifo_iarg_120_empty_n(ap_fifo_iarg_120_empty_n),
        .ap_fifo_iarg_120_dout(ap_fifo_iarg_120_dout),
        .ap_fifo_iarg_120_read(ap_fifo_iarg_120_read),
        .s_axis_fifo_121_tlast(s_axis_fifo_121_tlast),
        .s_axis_fifo_121_tvalid(s_axis_fifo_121_tvalid),
        .s_axis_fifo_121_tkeep(s_axis_fifo_121_tkeep),
        .s_axis_fifo_121_tstrb(s_axis_fifo_121_tstrb),
        .s_axis_fifo_121_tdata(s_axis_fifo_121_tdata),
        .s_axis_fifo_121_tready(s_axis_fifo_121_tready),
        .ap_fifo_iarg_121_empty_n(ap_fifo_iarg_121_empty_n),
        .ap_fifo_iarg_121_dout(ap_fifo_iarg_121_dout),
        .ap_fifo_iarg_121_read(ap_fifo_iarg_121_read),
        .s_axis_fifo_122_tlast(s_axis_fifo_122_tlast),
        .s_axis_fifo_122_tvalid(s_axis_fifo_122_tvalid),
        .s_axis_fifo_122_tkeep(s_axis_fifo_122_tkeep),
        .s_axis_fifo_122_tstrb(s_axis_fifo_122_tstrb),
        .s_axis_fifo_122_tdata(s_axis_fifo_122_tdata),
        .s_axis_fifo_122_tready(s_axis_fifo_122_tready),
        .ap_fifo_iarg_122_empty_n(ap_fifo_iarg_122_empty_n),
        .ap_fifo_iarg_122_dout(ap_fifo_iarg_122_dout),
        .ap_fifo_iarg_122_read(ap_fifo_iarg_122_read),
        .s_axis_fifo_123_tlast(s_axis_fifo_123_tlast),
        .s_axis_fifo_123_tvalid(s_axis_fifo_123_tvalid),
        .s_axis_fifo_123_tkeep(s_axis_fifo_123_tkeep),
        .s_axis_fifo_123_tstrb(s_axis_fifo_123_tstrb),
        .s_axis_fifo_123_tdata(s_axis_fifo_123_tdata),
        .s_axis_fifo_123_tready(s_axis_fifo_123_tready),
        .ap_fifo_iarg_123_empty_n(ap_fifo_iarg_123_empty_n),
        .ap_fifo_iarg_123_dout(ap_fifo_iarg_123_dout),
        .ap_fifo_iarg_123_read(ap_fifo_iarg_123_read),
        .s_axis_fifo_124_tlast(s_axis_fifo_124_tlast),
        .s_axis_fifo_124_tvalid(s_axis_fifo_124_tvalid),
        .s_axis_fifo_124_tkeep(s_axis_fifo_124_tkeep),
        .s_axis_fifo_124_tstrb(s_axis_fifo_124_tstrb),
        .s_axis_fifo_124_tdata(s_axis_fifo_124_tdata),
        .s_axis_fifo_124_tready(s_axis_fifo_124_tready),
        .ap_fifo_iarg_124_empty_n(ap_fifo_iarg_124_empty_n),
        .ap_fifo_iarg_124_dout(ap_fifo_iarg_124_dout),
        .ap_fifo_iarg_124_read(ap_fifo_iarg_124_read),
        .s_axis_fifo_125_tlast(s_axis_fifo_125_tlast),
        .s_axis_fifo_125_tvalid(s_axis_fifo_125_tvalid),
        .s_axis_fifo_125_tkeep(s_axis_fifo_125_tkeep),
        .s_axis_fifo_125_tstrb(s_axis_fifo_125_tstrb),
        .s_axis_fifo_125_tdata(s_axis_fifo_125_tdata),
        .s_axis_fifo_125_tready(s_axis_fifo_125_tready),
        .ap_fifo_iarg_125_empty_n(ap_fifo_iarg_125_empty_n),
        .ap_fifo_iarg_125_dout(ap_fifo_iarg_125_dout),
        .ap_fifo_iarg_125_read(ap_fifo_iarg_125_read),
        .s_axis_fifo_126_tlast(s_axis_fifo_126_tlast),
        .s_axis_fifo_126_tvalid(s_axis_fifo_126_tvalid),
        .s_axis_fifo_126_tkeep(s_axis_fifo_126_tkeep),
        .s_axis_fifo_126_tstrb(s_axis_fifo_126_tstrb),
        .s_axis_fifo_126_tdata(s_axis_fifo_126_tdata),
        .s_axis_fifo_126_tready(s_axis_fifo_126_tready),
        .ap_fifo_iarg_126_empty_n(ap_fifo_iarg_126_empty_n),
        .ap_fifo_iarg_126_dout(ap_fifo_iarg_126_dout),
        .ap_fifo_iarg_126_read(ap_fifo_iarg_126_read),
        .s_axis_fifo_127_tlast(s_axis_fifo_127_tlast),
        .s_axis_fifo_127_tvalid(s_axis_fifo_127_tvalid),
        .s_axis_fifo_127_tkeep(s_axis_fifo_127_tkeep),
        .s_axis_fifo_127_tstrb(s_axis_fifo_127_tstrb),
        .s_axis_fifo_127_tdata(s_axis_fifo_127_tdata),
        .s_axis_fifo_127_tready(s_axis_fifo_127_tready),
        .ap_fifo_iarg_127_empty_n(ap_fifo_iarg_127_empty_n),
        .ap_fifo_iarg_127_dout(ap_fifo_iarg_127_dout),
        .ap_fifo_iarg_127_read(ap_fifo_iarg_127_read)
    );
        
    out_fifo_args #(
        .C_NUM_OUTPUT_FIFOs(C_NUM_OUTPUT_FIFOs),
        .C_OUTPUT_FIFO_0_WIDTH(C_OUTPUT_FIFO_0_WIDTH),
        .C_OUTPUT_FIFO_1_WIDTH(C_OUTPUT_FIFO_1_WIDTH),
        .C_OUTPUT_FIFO_2_WIDTH(C_OUTPUT_FIFO_2_WIDTH),
        .C_OUTPUT_FIFO_3_WIDTH(C_OUTPUT_FIFO_3_WIDTH),
        .C_OUTPUT_FIFO_4_WIDTH(C_OUTPUT_FIFO_4_WIDTH),
        .C_OUTPUT_FIFO_5_WIDTH(C_OUTPUT_FIFO_5_WIDTH),
        .C_OUTPUT_FIFO_6_WIDTH(C_OUTPUT_FIFO_6_WIDTH),
        .C_OUTPUT_FIFO_7_WIDTH(C_OUTPUT_FIFO_7_WIDTH),
        .C_OUTPUT_FIFO_8_WIDTH(C_OUTPUT_FIFO_8_WIDTH),
        .C_OUTPUT_FIFO_9_WIDTH(C_OUTPUT_FIFO_9_WIDTH),
        .C_OUTPUT_FIFO_10_WIDTH(C_OUTPUT_FIFO_10_WIDTH),
        .C_OUTPUT_FIFO_11_WIDTH(C_OUTPUT_FIFO_11_WIDTH),
        .C_OUTPUT_FIFO_12_WIDTH(C_OUTPUT_FIFO_12_WIDTH),
        .C_OUTPUT_FIFO_13_WIDTH(C_OUTPUT_FIFO_13_WIDTH),
        .C_OUTPUT_FIFO_14_WIDTH(C_OUTPUT_FIFO_14_WIDTH),
        .C_OUTPUT_FIFO_15_WIDTH(C_OUTPUT_FIFO_15_WIDTH),
        .C_OUTPUT_FIFO_16_WIDTH(C_OUTPUT_FIFO_16_WIDTH),
        .C_OUTPUT_FIFO_17_WIDTH(C_OUTPUT_FIFO_17_WIDTH),
        .C_OUTPUT_FIFO_18_WIDTH(C_OUTPUT_FIFO_18_WIDTH),
        .C_OUTPUT_FIFO_19_WIDTH(C_OUTPUT_FIFO_19_WIDTH),
        .C_OUTPUT_FIFO_20_WIDTH(C_OUTPUT_FIFO_20_WIDTH),
        .C_OUTPUT_FIFO_21_WIDTH(C_OUTPUT_FIFO_21_WIDTH),
        .C_OUTPUT_FIFO_22_WIDTH(C_OUTPUT_FIFO_22_WIDTH),
        .C_OUTPUT_FIFO_23_WIDTH(C_OUTPUT_FIFO_23_WIDTH),
        .C_OUTPUT_FIFO_24_WIDTH(C_OUTPUT_FIFO_24_WIDTH),
        .C_OUTPUT_FIFO_25_WIDTH(C_OUTPUT_FIFO_25_WIDTH),
        .C_OUTPUT_FIFO_26_WIDTH(C_OUTPUT_FIFO_26_WIDTH),
        .C_OUTPUT_FIFO_27_WIDTH(C_OUTPUT_FIFO_27_WIDTH),
        .C_OUTPUT_FIFO_28_WIDTH(C_OUTPUT_FIFO_28_WIDTH),
        .C_OUTPUT_FIFO_29_WIDTH(C_OUTPUT_FIFO_29_WIDTH),
        .C_OUTPUT_FIFO_30_WIDTH(C_OUTPUT_FIFO_30_WIDTH),
        .C_OUTPUT_FIFO_31_WIDTH(C_OUTPUT_FIFO_31_WIDTH),
        .C_OUTPUT_FIFO_32_WIDTH(C_OUTPUT_FIFO_32_WIDTH),
        .C_OUTPUT_FIFO_33_WIDTH(C_OUTPUT_FIFO_33_WIDTH),
        .C_OUTPUT_FIFO_34_WIDTH(C_OUTPUT_FIFO_34_WIDTH),
        .C_OUTPUT_FIFO_35_WIDTH(C_OUTPUT_FIFO_35_WIDTH),
        .C_OUTPUT_FIFO_36_WIDTH(C_OUTPUT_FIFO_36_WIDTH),
        .C_OUTPUT_FIFO_37_WIDTH(C_OUTPUT_FIFO_37_WIDTH),
        .C_OUTPUT_FIFO_38_WIDTH(C_OUTPUT_FIFO_38_WIDTH),
        .C_OUTPUT_FIFO_39_WIDTH(C_OUTPUT_FIFO_39_WIDTH),
        .C_OUTPUT_FIFO_40_WIDTH(C_OUTPUT_FIFO_40_WIDTH),
        .C_OUTPUT_FIFO_41_WIDTH(C_OUTPUT_FIFO_41_WIDTH),
        .C_OUTPUT_FIFO_42_WIDTH(C_OUTPUT_FIFO_42_WIDTH),
        .C_OUTPUT_FIFO_43_WIDTH(C_OUTPUT_FIFO_43_WIDTH),
        .C_OUTPUT_FIFO_44_WIDTH(C_OUTPUT_FIFO_44_WIDTH),
        .C_OUTPUT_FIFO_45_WIDTH(C_OUTPUT_FIFO_45_WIDTH),
        .C_OUTPUT_FIFO_46_WIDTH(C_OUTPUT_FIFO_46_WIDTH),
        .C_OUTPUT_FIFO_47_WIDTH(C_OUTPUT_FIFO_47_WIDTH),
        .C_OUTPUT_FIFO_48_WIDTH(C_OUTPUT_FIFO_48_WIDTH),
        .C_OUTPUT_FIFO_49_WIDTH(C_OUTPUT_FIFO_49_WIDTH),
        .C_OUTPUT_FIFO_50_WIDTH(C_OUTPUT_FIFO_50_WIDTH),
        .C_OUTPUT_FIFO_51_WIDTH(C_OUTPUT_FIFO_51_WIDTH),
        .C_OUTPUT_FIFO_52_WIDTH(C_OUTPUT_FIFO_52_WIDTH),
        .C_OUTPUT_FIFO_53_WIDTH(C_OUTPUT_FIFO_53_WIDTH),
        .C_OUTPUT_FIFO_54_WIDTH(C_OUTPUT_FIFO_54_WIDTH),
        .C_OUTPUT_FIFO_55_WIDTH(C_OUTPUT_FIFO_55_WIDTH),
        .C_OUTPUT_FIFO_56_WIDTH(C_OUTPUT_FIFO_56_WIDTH),
        .C_OUTPUT_FIFO_57_WIDTH(C_OUTPUT_FIFO_57_WIDTH),
        .C_OUTPUT_FIFO_58_WIDTH(C_OUTPUT_FIFO_58_WIDTH),
        .C_OUTPUT_FIFO_59_WIDTH(C_OUTPUT_FIFO_59_WIDTH),
        .C_OUTPUT_FIFO_60_WIDTH(C_OUTPUT_FIFO_60_WIDTH),
        .C_OUTPUT_FIFO_61_WIDTH(C_OUTPUT_FIFO_61_WIDTH),
        .C_OUTPUT_FIFO_62_WIDTH(C_OUTPUT_FIFO_62_WIDTH),
        .C_OUTPUT_FIFO_63_WIDTH(C_OUTPUT_FIFO_63_WIDTH),
        .C_OUTPUT_FIFO_64_WIDTH(C_OUTPUT_FIFO_64_WIDTH),
        .C_OUTPUT_FIFO_65_WIDTH(C_OUTPUT_FIFO_65_WIDTH),
        .C_OUTPUT_FIFO_66_WIDTH(C_OUTPUT_FIFO_66_WIDTH),
        .C_OUTPUT_FIFO_67_WIDTH(C_OUTPUT_FIFO_67_WIDTH),
        .C_OUTPUT_FIFO_68_WIDTH(C_OUTPUT_FIFO_68_WIDTH),
        .C_OUTPUT_FIFO_69_WIDTH(C_OUTPUT_FIFO_69_WIDTH),
        .C_OUTPUT_FIFO_70_WIDTH(C_OUTPUT_FIFO_70_WIDTH),
        .C_OUTPUT_FIFO_71_WIDTH(C_OUTPUT_FIFO_71_WIDTH),
        .C_OUTPUT_FIFO_72_WIDTH(C_OUTPUT_FIFO_72_WIDTH),
        .C_OUTPUT_FIFO_73_WIDTH(C_OUTPUT_FIFO_73_WIDTH),
        .C_OUTPUT_FIFO_74_WIDTH(C_OUTPUT_FIFO_74_WIDTH),
        .C_OUTPUT_FIFO_75_WIDTH(C_OUTPUT_FIFO_75_WIDTH),
        .C_OUTPUT_FIFO_76_WIDTH(C_OUTPUT_FIFO_76_WIDTH),
        .C_OUTPUT_FIFO_77_WIDTH(C_OUTPUT_FIFO_77_WIDTH),
        .C_OUTPUT_FIFO_78_WIDTH(C_OUTPUT_FIFO_78_WIDTH),
        .C_OUTPUT_FIFO_79_WIDTH(C_OUTPUT_FIFO_79_WIDTH),
        .C_OUTPUT_FIFO_80_WIDTH(C_OUTPUT_FIFO_80_WIDTH),
        .C_OUTPUT_FIFO_81_WIDTH(C_OUTPUT_FIFO_81_WIDTH),
        .C_OUTPUT_FIFO_82_WIDTH(C_OUTPUT_FIFO_82_WIDTH),
        .C_OUTPUT_FIFO_83_WIDTH(C_OUTPUT_FIFO_83_WIDTH),
        .C_OUTPUT_FIFO_84_WIDTH(C_OUTPUT_FIFO_84_WIDTH),
        .C_OUTPUT_FIFO_85_WIDTH(C_OUTPUT_FIFO_85_WIDTH),
        .C_OUTPUT_FIFO_86_WIDTH(C_OUTPUT_FIFO_86_WIDTH),
        .C_OUTPUT_FIFO_87_WIDTH(C_OUTPUT_FIFO_87_WIDTH),
        .C_OUTPUT_FIFO_88_WIDTH(C_OUTPUT_FIFO_88_WIDTH),
        .C_OUTPUT_FIFO_89_WIDTH(C_OUTPUT_FIFO_89_WIDTH),
        .C_OUTPUT_FIFO_90_WIDTH(C_OUTPUT_FIFO_90_WIDTH),
        .C_OUTPUT_FIFO_91_WIDTH(C_OUTPUT_FIFO_91_WIDTH),
        .C_OUTPUT_FIFO_92_WIDTH(C_OUTPUT_FIFO_92_WIDTH),
        .C_OUTPUT_FIFO_93_WIDTH(C_OUTPUT_FIFO_93_WIDTH),
        .C_OUTPUT_FIFO_94_WIDTH(C_OUTPUT_FIFO_94_WIDTH),
        .C_OUTPUT_FIFO_95_WIDTH(C_OUTPUT_FIFO_95_WIDTH),
        .C_OUTPUT_FIFO_96_WIDTH(C_OUTPUT_FIFO_96_WIDTH),
        .C_OUTPUT_FIFO_97_WIDTH(C_OUTPUT_FIFO_97_WIDTH),
        .C_OUTPUT_FIFO_98_WIDTH(C_OUTPUT_FIFO_98_WIDTH),
        .C_OUTPUT_FIFO_99_WIDTH(C_OUTPUT_FIFO_99_WIDTH),
        .C_OUTPUT_FIFO_100_WIDTH(C_OUTPUT_FIFO_100_WIDTH),
        .C_OUTPUT_FIFO_101_WIDTH(C_OUTPUT_FIFO_101_WIDTH),
        .C_OUTPUT_FIFO_102_WIDTH(C_OUTPUT_FIFO_102_WIDTH),
        .C_OUTPUT_FIFO_103_WIDTH(C_OUTPUT_FIFO_103_WIDTH),
        .C_OUTPUT_FIFO_104_WIDTH(C_OUTPUT_FIFO_104_WIDTH),
        .C_OUTPUT_FIFO_105_WIDTH(C_OUTPUT_FIFO_105_WIDTH),
        .C_OUTPUT_FIFO_106_WIDTH(C_OUTPUT_FIFO_106_WIDTH),
        .C_OUTPUT_FIFO_107_WIDTH(C_OUTPUT_FIFO_107_WIDTH),
        .C_OUTPUT_FIFO_108_WIDTH(C_OUTPUT_FIFO_108_WIDTH),
        .C_OUTPUT_FIFO_109_WIDTH(C_OUTPUT_FIFO_109_WIDTH),
        .C_OUTPUT_FIFO_110_WIDTH(C_OUTPUT_FIFO_110_WIDTH),
        .C_OUTPUT_FIFO_111_WIDTH(C_OUTPUT_FIFO_111_WIDTH),
        .C_OUTPUT_FIFO_112_WIDTH(C_OUTPUT_FIFO_112_WIDTH),
        .C_OUTPUT_FIFO_113_WIDTH(C_OUTPUT_FIFO_113_WIDTH),
        .C_OUTPUT_FIFO_114_WIDTH(C_OUTPUT_FIFO_114_WIDTH),
        .C_OUTPUT_FIFO_115_WIDTH(C_OUTPUT_FIFO_115_WIDTH),
        .C_OUTPUT_FIFO_116_WIDTH(C_OUTPUT_FIFO_116_WIDTH),
        .C_OUTPUT_FIFO_117_WIDTH(C_OUTPUT_FIFO_117_WIDTH),
        .C_OUTPUT_FIFO_118_WIDTH(C_OUTPUT_FIFO_118_WIDTH),
        .C_OUTPUT_FIFO_119_WIDTH(C_OUTPUT_FIFO_119_WIDTH),
        .C_OUTPUT_FIFO_120_WIDTH(C_OUTPUT_FIFO_120_WIDTH),
        .C_OUTPUT_FIFO_121_WIDTH(C_OUTPUT_FIFO_121_WIDTH),
        .C_OUTPUT_FIFO_122_WIDTH(C_OUTPUT_FIFO_122_WIDTH),
        .C_OUTPUT_FIFO_123_WIDTH(C_OUTPUT_FIFO_123_WIDTH),
        .C_OUTPUT_FIFO_124_WIDTH(C_OUTPUT_FIFO_124_WIDTH),
        .C_OUTPUT_FIFO_125_WIDTH(C_OUTPUT_FIFO_125_WIDTH),
        .C_OUTPUT_FIFO_126_WIDTH(C_OUTPUT_FIFO_126_WIDTH),
        .C_OUTPUT_FIFO_127_WIDTH(C_OUTPUT_FIFO_127_WIDTH),
        .C_OUTPUT_FIFO_0_DEPTH(C_OUTPUT_FIFO_0_DEPTH),
        .C_OUTPUT_FIFO_1_DEPTH(C_OUTPUT_FIFO_1_DEPTH),
        .C_OUTPUT_FIFO_2_DEPTH(C_OUTPUT_FIFO_2_DEPTH),
        .C_OUTPUT_FIFO_3_DEPTH(C_OUTPUT_FIFO_3_DEPTH),
        .C_OUTPUT_FIFO_4_DEPTH(C_OUTPUT_FIFO_4_DEPTH),
        .C_OUTPUT_FIFO_5_DEPTH(C_OUTPUT_FIFO_5_DEPTH),
        .C_OUTPUT_FIFO_6_DEPTH(C_OUTPUT_FIFO_6_DEPTH),
        .C_OUTPUT_FIFO_7_DEPTH(C_OUTPUT_FIFO_7_DEPTH),
        .C_OUTPUT_FIFO_8_DEPTH(C_OUTPUT_FIFO_8_DEPTH),
        .C_OUTPUT_FIFO_9_DEPTH(C_OUTPUT_FIFO_9_DEPTH),
        .C_OUTPUT_FIFO_10_DEPTH(C_OUTPUT_FIFO_10_DEPTH),
        .C_OUTPUT_FIFO_11_DEPTH(C_OUTPUT_FIFO_11_DEPTH),
        .C_OUTPUT_FIFO_12_DEPTH(C_OUTPUT_FIFO_12_DEPTH),
        .C_OUTPUT_FIFO_13_DEPTH(C_OUTPUT_FIFO_13_DEPTH),
        .C_OUTPUT_FIFO_14_DEPTH(C_OUTPUT_FIFO_14_DEPTH),
        .C_OUTPUT_FIFO_15_DEPTH(C_OUTPUT_FIFO_15_DEPTH),
        .C_OUTPUT_FIFO_16_DEPTH(C_OUTPUT_FIFO_16_DEPTH),
        .C_OUTPUT_FIFO_17_DEPTH(C_OUTPUT_FIFO_17_DEPTH),
        .C_OUTPUT_FIFO_18_DEPTH(C_OUTPUT_FIFO_18_DEPTH),
        .C_OUTPUT_FIFO_19_DEPTH(C_OUTPUT_FIFO_19_DEPTH),
        .C_OUTPUT_FIFO_20_DEPTH(C_OUTPUT_FIFO_20_DEPTH),
        .C_OUTPUT_FIFO_21_DEPTH(C_OUTPUT_FIFO_21_DEPTH),
        .C_OUTPUT_FIFO_22_DEPTH(C_OUTPUT_FIFO_22_DEPTH),
        .C_OUTPUT_FIFO_23_DEPTH(C_OUTPUT_FIFO_23_DEPTH),
        .C_OUTPUT_FIFO_24_DEPTH(C_OUTPUT_FIFO_24_DEPTH),
        .C_OUTPUT_FIFO_25_DEPTH(C_OUTPUT_FIFO_25_DEPTH),
        .C_OUTPUT_FIFO_26_DEPTH(C_OUTPUT_FIFO_26_DEPTH),
        .C_OUTPUT_FIFO_27_DEPTH(C_OUTPUT_FIFO_27_DEPTH),
        .C_OUTPUT_FIFO_28_DEPTH(C_OUTPUT_FIFO_28_DEPTH),
        .C_OUTPUT_FIFO_29_DEPTH(C_OUTPUT_FIFO_29_DEPTH),
        .C_OUTPUT_FIFO_30_DEPTH(C_OUTPUT_FIFO_30_DEPTH),
        .C_OUTPUT_FIFO_31_DEPTH(C_OUTPUT_FIFO_31_DEPTH),
        .C_OUTPUT_FIFO_32_DEPTH(C_OUTPUT_FIFO_32_DEPTH),
        .C_OUTPUT_FIFO_33_DEPTH(C_OUTPUT_FIFO_33_DEPTH),
        .C_OUTPUT_FIFO_34_DEPTH(C_OUTPUT_FIFO_34_DEPTH),
        .C_OUTPUT_FIFO_35_DEPTH(C_OUTPUT_FIFO_35_DEPTH),
        .C_OUTPUT_FIFO_36_DEPTH(C_OUTPUT_FIFO_36_DEPTH),
        .C_OUTPUT_FIFO_37_DEPTH(C_OUTPUT_FIFO_37_DEPTH),
        .C_OUTPUT_FIFO_38_DEPTH(C_OUTPUT_FIFO_38_DEPTH),
        .C_OUTPUT_FIFO_39_DEPTH(C_OUTPUT_FIFO_39_DEPTH),
        .C_OUTPUT_FIFO_40_DEPTH(C_OUTPUT_FIFO_40_DEPTH),
        .C_OUTPUT_FIFO_41_DEPTH(C_OUTPUT_FIFO_41_DEPTH),
        .C_OUTPUT_FIFO_42_DEPTH(C_OUTPUT_FIFO_42_DEPTH),
        .C_OUTPUT_FIFO_43_DEPTH(C_OUTPUT_FIFO_43_DEPTH),
        .C_OUTPUT_FIFO_44_DEPTH(C_OUTPUT_FIFO_44_DEPTH),
        .C_OUTPUT_FIFO_45_DEPTH(C_OUTPUT_FIFO_45_DEPTH),
        .C_OUTPUT_FIFO_46_DEPTH(C_OUTPUT_FIFO_46_DEPTH),
        .C_OUTPUT_FIFO_47_DEPTH(C_OUTPUT_FIFO_47_DEPTH),
        .C_OUTPUT_FIFO_48_DEPTH(C_OUTPUT_FIFO_48_DEPTH),
        .C_OUTPUT_FIFO_49_DEPTH(C_OUTPUT_FIFO_49_DEPTH),
        .C_OUTPUT_FIFO_50_DEPTH(C_OUTPUT_FIFO_50_DEPTH),
        .C_OUTPUT_FIFO_51_DEPTH(C_OUTPUT_FIFO_51_DEPTH),
        .C_OUTPUT_FIFO_52_DEPTH(C_OUTPUT_FIFO_52_DEPTH),
        .C_OUTPUT_FIFO_53_DEPTH(C_OUTPUT_FIFO_53_DEPTH),
        .C_OUTPUT_FIFO_54_DEPTH(C_OUTPUT_FIFO_54_DEPTH),
        .C_OUTPUT_FIFO_55_DEPTH(C_OUTPUT_FIFO_55_DEPTH),
        .C_OUTPUT_FIFO_56_DEPTH(C_OUTPUT_FIFO_56_DEPTH),
        .C_OUTPUT_FIFO_57_DEPTH(C_OUTPUT_FIFO_57_DEPTH),
        .C_OUTPUT_FIFO_58_DEPTH(C_OUTPUT_FIFO_58_DEPTH),
        .C_OUTPUT_FIFO_59_DEPTH(C_OUTPUT_FIFO_59_DEPTH),
        .C_OUTPUT_FIFO_60_DEPTH(C_OUTPUT_FIFO_60_DEPTH),
        .C_OUTPUT_FIFO_61_DEPTH(C_OUTPUT_FIFO_61_DEPTH),
        .C_OUTPUT_FIFO_62_DEPTH(C_OUTPUT_FIFO_62_DEPTH),
        .C_OUTPUT_FIFO_63_DEPTH(C_OUTPUT_FIFO_63_DEPTH),
        .C_OUTPUT_FIFO_64_DEPTH(C_OUTPUT_FIFO_64_DEPTH),
        .C_OUTPUT_FIFO_65_DEPTH(C_OUTPUT_FIFO_65_DEPTH),
        .C_OUTPUT_FIFO_66_DEPTH(C_OUTPUT_FIFO_66_DEPTH),
        .C_OUTPUT_FIFO_67_DEPTH(C_OUTPUT_FIFO_67_DEPTH),
        .C_OUTPUT_FIFO_68_DEPTH(C_OUTPUT_FIFO_68_DEPTH),
        .C_OUTPUT_FIFO_69_DEPTH(C_OUTPUT_FIFO_69_DEPTH),
        .C_OUTPUT_FIFO_70_DEPTH(C_OUTPUT_FIFO_70_DEPTH),
        .C_OUTPUT_FIFO_71_DEPTH(C_OUTPUT_FIFO_71_DEPTH),
        .C_OUTPUT_FIFO_72_DEPTH(C_OUTPUT_FIFO_72_DEPTH),
        .C_OUTPUT_FIFO_73_DEPTH(C_OUTPUT_FIFO_73_DEPTH),
        .C_OUTPUT_FIFO_74_DEPTH(C_OUTPUT_FIFO_74_DEPTH),
        .C_OUTPUT_FIFO_75_DEPTH(C_OUTPUT_FIFO_75_DEPTH),
        .C_OUTPUT_FIFO_76_DEPTH(C_OUTPUT_FIFO_76_DEPTH),
        .C_OUTPUT_FIFO_77_DEPTH(C_OUTPUT_FIFO_77_DEPTH),
        .C_OUTPUT_FIFO_78_DEPTH(C_OUTPUT_FIFO_78_DEPTH),
        .C_OUTPUT_FIFO_79_DEPTH(C_OUTPUT_FIFO_79_DEPTH),
        .C_OUTPUT_FIFO_80_DEPTH(C_OUTPUT_FIFO_80_DEPTH),
        .C_OUTPUT_FIFO_81_DEPTH(C_OUTPUT_FIFO_81_DEPTH),
        .C_OUTPUT_FIFO_82_DEPTH(C_OUTPUT_FIFO_82_DEPTH),
        .C_OUTPUT_FIFO_83_DEPTH(C_OUTPUT_FIFO_83_DEPTH),
        .C_OUTPUT_FIFO_84_DEPTH(C_OUTPUT_FIFO_84_DEPTH),
        .C_OUTPUT_FIFO_85_DEPTH(C_OUTPUT_FIFO_85_DEPTH),
        .C_OUTPUT_FIFO_86_DEPTH(C_OUTPUT_FIFO_86_DEPTH),
        .C_OUTPUT_FIFO_87_DEPTH(C_OUTPUT_FIFO_87_DEPTH),
        .C_OUTPUT_FIFO_88_DEPTH(C_OUTPUT_FIFO_88_DEPTH),
        .C_OUTPUT_FIFO_89_DEPTH(C_OUTPUT_FIFO_89_DEPTH),
        .C_OUTPUT_FIFO_90_DEPTH(C_OUTPUT_FIFO_90_DEPTH),
        .C_OUTPUT_FIFO_91_DEPTH(C_OUTPUT_FIFO_91_DEPTH),
        .C_OUTPUT_FIFO_92_DEPTH(C_OUTPUT_FIFO_92_DEPTH),
        .C_OUTPUT_FIFO_93_DEPTH(C_OUTPUT_FIFO_93_DEPTH),
        .C_OUTPUT_FIFO_94_DEPTH(C_OUTPUT_FIFO_94_DEPTH),
        .C_OUTPUT_FIFO_95_DEPTH(C_OUTPUT_FIFO_95_DEPTH),
        .C_OUTPUT_FIFO_96_DEPTH(C_OUTPUT_FIFO_96_DEPTH),
        .C_OUTPUT_FIFO_97_DEPTH(C_OUTPUT_FIFO_97_DEPTH),
        .C_OUTPUT_FIFO_98_DEPTH(C_OUTPUT_FIFO_98_DEPTH),
        .C_OUTPUT_FIFO_99_DEPTH(C_OUTPUT_FIFO_99_DEPTH),
        .C_OUTPUT_FIFO_100_DEPTH(C_OUTPUT_FIFO_100_DEPTH),
        .C_OUTPUT_FIFO_101_DEPTH(C_OUTPUT_FIFO_101_DEPTH),
        .C_OUTPUT_FIFO_102_DEPTH(C_OUTPUT_FIFO_102_DEPTH),
        .C_OUTPUT_FIFO_103_DEPTH(C_OUTPUT_FIFO_103_DEPTH),
        .C_OUTPUT_FIFO_104_DEPTH(C_OUTPUT_FIFO_104_DEPTH),
        .C_OUTPUT_FIFO_105_DEPTH(C_OUTPUT_FIFO_105_DEPTH),
        .C_OUTPUT_FIFO_106_DEPTH(C_OUTPUT_FIFO_106_DEPTH),
        .C_OUTPUT_FIFO_107_DEPTH(C_OUTPUT_FIFO_107_DEPTH),
        .C_OUTPUT_FIFO_108_DEPTH(C_OUTPUT_FIFO_108_DEPTH),
        .C_OUTPUT_FIFO_109_DEPTH(C_OUTPUT_FIFO_109_DEPTH),
        .C_OUTPUT_FIFO_110_DEPTH(C_OUTPUT_FIFO_110_DEPTH),
        .C_OUTPUT_FIFO_111_DEPTH(C_OUTPUT_FIFO_111_DEPTH),
        .C_OUTPUT_FIFO_112_DEPTH(C_OUTPUT_FIFO_112_DEPTH),
        .C_OUTPUT_FIFO_113_DEPTH(C_OUTPUT_FIFO_113_DEPTH),
        .C_OUTPUT_FIFO_114_DEPTH(C_OUTPUT_FIFO_114_DEPTH),
        .C_OUTPUT_FIFO_115_DEPTH(C_OUTPUT_FIFO_115_DEPTH),
        .C_OUTPUT_FIFO_116_DEPTH(C_OUTPUT_FIFO_116_DEPTH),
        .C_OUTPUT_FIFO_117_DEPTH(C_OUTPUT_FIFO_117_DEPTH),
        .C_OUTPUT_FIFO_118_DEPTH(C_OUTPUT_FIFO_118_DEPTH),
        .C_OUTPUT_FIFO_119_DEPTH(C_OUTPUT_FIFO_119_DEPTH),
        .C_OUTPUT_FIFO_120_DEPTH(C_OUTPUT_FIFO_120_DEPTH),
        .C_OUTPUT_FIFO_121_DEPTH(C_OUTPUT_FIFO_121_DEPTH),
        .C_OUTPUT_FIFO_122_DEPTH(C_OUTPUT_FIFO_122_DEPTH),
        .C_OUTPUT_FIFO_123_DEPTH(C_OUTPUT_FIFO_123_DEPTH),
        .C_OUTPUT_FIFO_124_DEPTH(C_OUTPUT_FIFO_124_DEPTH),
        .C_OUTPUT_FIFO_125_DEPTH(C_OUTPUT_FIFO_125_DEPTH),
        .C_OUTPUT_FIFO_126_DEPTH(C_OUTPUT_FIFO_126_DEPTH),
        .C_OUTPUT_FIFO_127_DEPTH(C_OUTPUT_FIFO_127_DEPTH),
        .C_OUTPUT_FIFO_0_DMWIDTH(C_OUTPUT_FIFO_0_DMWIDTH),
        .C_OUTPUT_FIFO_1_DMWIDTH(C_OUTPUT_FIFO_1_DMWIDTH),
        .C_OUTPUT_FIFO_2_DMWIDTH(C_OUTPUT_FIFO_2_DMWIDTH),
        .C_OUTPUT_FIFO_3_DMWIDTH(C_OUTPUT_FIFO_3_DMWIDTH),
        .C_OUTPUT_FIFO_4_DMWIDTH(C_OUTPUT_FIFO_4_DMWIDTH),
        .C_OUTPUT_FIFO_5_DMWIDTH(C_OUTPUT_FIFO_5_DMWIDTH),
        .C_OUTPUT_FIFO_6_DMWIDTH(C_OUTPUT_FIFO_6_DMWIDTH),
        .C_OUTPUT_FIFO_7_DMWIDTH(C_OUTPUT_FIFO_7_DMWIDTH),
        .C_OUTPUT_FIFO_8_DMWIDTH(C_OUTPUT_FIFO_8_DMWIDTH),
        .C_OUTPUT_FIFO_9_DMWIDTH(C_OUTPUT_FIFO_9_DMWIDTH),
        .C_OUTPUT_FIFO_10_DMWIDTH(C_OUTPUT_FIFO_10_DMWIDTH),
        .C_OUTPUT_FIFO_11_DMWIDTH(C_OUTPUT_FIFO_11_DMWIDTH),
        .C_OUTPUT_FIFO_12_DMWIDTH(C_OUTPUT_FIFO_12_DMWIDTH),
        .C_OUTPUT_FIFO_13_DMWIDTH(C_OUTPUT_FIFO_13_DMWIDTH),
        .C_OUTPUT_FIFO_14_DMWIDTH(C_OUTPUT_FIFO_14_DMWIDTH),
        .C_OUTPUT_FIFO_15_DMWIDTH(C_OUTPUT_FIFO_15_DMWIDTH),
        .C_OUTPUT_FIFO_16_DMWIDTH(C_OUTPUT_FIFO_16_DMWIDTH),
        .C_OUTPUT_FIFO_17_DMWIDTH(C_OUTPUT_FIFO_17_DMWIDTH),
        .C_OUTPUT_FIFO_18_DMWIDTH(C_OUTPUT_FIFO_18_DMWIDTH),
        .C_OUTPUT_FIFO_19_DMWIDTH(C_OUTPUT_FIFO_19_DMWIDTH),
        .C_OUTPUT_FIFO_20_DMWIDTH(C_OUTPUT_FIFO_20_DMWIDTH),
        .C_OUTPUT_FIFO_21_DMWIDTH(C_OUTPUT_FIFO_21_DMWIDTH),
        .C_OUTPUT_FIFO_22_DMWIDTH(C_OUTPUT_FIFO_22_DMWIDTH),
        .C_OUTPUT_FIFO_23_DMWIDTH(C_OUTPUT_FIFO_23_DMWIDTH),
        .C_OUTPUT_FIFO_24_DMWIDTH(C_OUTPUT_FIFO_24_DMWIDTH),
        .C_OUTPUT_FIFO_25_DMWIDTH(C_OUTPUT_FIFO_25_DMWIDTH),
        .C_OUTPUT_FIFO_26_DMWIDTH(C_OUTPUT_FIFO_26_DMWIDTH),
        .C_OUTPUT_FIFO_27_DMWIDTH(C_OUTPUT_FIFO_27_DMWIDTH),
        .C_OUTPUT_FIFO_28_DMWIDTH(C_OUTPUT_FIFO_28_DMWIDTH),
        .C_OUTPUT_FIFO_29_DMWIDTH(C_OUTPUT_FIFO_29_DMWIDTH),
        .C_OUTPUT_FIFO_30_DMWIDTH(C_OUTPUT_FIFO_30_DMWIDTH),
        .C_OUTPUT_FIFO_31_DMWIDTH(C_OUTPUT_FIFO_31_DMWIDTH),
        .C_OUTPUT_FIFO_32_DMWIDTH(C_OUTPUT_FIFO_32_DMWIDTH),
        .C_OUTPUT_FIFO_33_DMWIDTH(C_OUTPUT_FIFO_33_DMWIDTH),
        .C_OUTPUT_FIFO_34_DMWIDTH(C_OUTPUT_FIFO_34_DMWIDTH),
        .C_OUTPUT_FIFO_35_DMWIDTH(C_OUTPUT_FIFO_35_DMWIDTH),
        .C_OUTPUT_FIFO_36_DMWIDTH(C_OUTPUT_FIFO_36_DMWIDTH),
        .C_OUTPUT_FIFO_37_DMWIDTH(C_OUTPUT_FIFO_37_DMWIDTH),
        .C_OUTPUT_FIFO_38_DMWIDTH(C_OUTPUT_FIFO_38_DMWIDTH),
        .C_OUTPUT_FIFO_39_DMWIDTH(C_OUTPUT_FIFO_39_DMWIDTH),
        .C_OUTPUT_FIFO_40_DMWIDTH(C_OUTPUT_FIFO_40_DMWIDTH),
        .C_OUTPUT_FIFO_41_DMWIDTH(C_OUTPUT_FIFO_41_DMWIDTH),
        .C_OUTPUT_FIFO_42_DMWIDTH(C_OUTPUT_FIFO_42_DMWIDTH),
        .C_OUTPUT_FIFO_43_DMWIDTH(C_OUTPUT_FIFO_43_DMWIDTH),
        .C_OUTPUT_FIFO_44_DMWIDTH(C_OUTPUT_FIFO_44_DMWIDTH),
        .C_OUTPUT_FIFO_45_DMWIDTH(C_OUTPUT_FIFO_45_DMWIDTH),
        .C_OUTPUT_FIFO_46_DMWIDTH(C_OUTPUT_FIFO_46_DMWIDTH),
        .C_OUTPUT_FIFO_47_DMWIDTH(C_OUTPUT_FIFO_47_DMWIDTH),
        .C_OUTPUT_FIFO_48_DMWIDTH(C_OUTPUT_FIFO_48_DMWIDTH),
        .C_OUTPUT_FIFO_49_DMWIDTH(C_OUTPUT_FIFO_49_DMWIDTH),
        .C_OUTPUT_FIFO_50_DMWIDTH(C_OUTPUT_FIFO_50_DMWIDTH),
        .C_OUTPUT_FIFO_51_DMWIDTH(C_OUTPUT_FIFO_51_DMWIDTH),
        .C_OUTPUT_FIFO_52_DMWIDTH(C_OUTPUT_FIFO_52_DMWIDTH),
        .C_OUTPUT_FIFO_53_DMWIDTH(C_OUTPUT_FIFO_53_DMWIDTH),
        .C_OUTPUT_FIFO_54_DMWIDTH(C_OUTPUT_FIFO_54_DMWIDTH),
        .C_OUTPUT_FIFO_55_DMWIDTH(C_OUTPUT_FIFO_55_DMWIDTH),
        .C_OUTPUT_FIFO_56_DMWIDTH(C_OUTPUT_FIFO_56_DMWIDTH),
        .C_OUTPUT_FIFO_57_DMWIDTH(C_OUTPUT_FIFO_57_DMWIDTH),
        .C_OUTPUT_FIFO_58_DMWIDTH(C_OUTPUT_FIFO_58_DMWIDTH),
        .C_OUTPUT_FIFO_59_DMWIDTH(C_OUTPUT_FIFO_59_DMWIDTH),
        .C_OUTPUT_FIFO_60_DMWIDTH(C_OUTPUT_FIFO_60_DMWIDTH),
        .C_OUTPUT_FIFO_61_DMWIDTH(C_OUTPUT_FIFO_61_DMWIDTH),
        .C_OUTPUT_FIFO_62_DMWIDTH(C_OUTPUT_FIFO_62_DMWIDTH),
        .C_OUTPUT_FIFO_63_DMWIDTH(C_OUTPUT_FIFO_63_DMWIDTH),
        .C_OUTPUT_FIFO_64_DMWIDTH(C_OUTPUT_FIFO_64_DMWIDTH),
        .C_OUTPUT_FIFO_65_DMWIDTH(C_OUTPUT_FIFO_65_DMWIDTH),
        .C_OUTPUT_FIFO_66_DMWIDTH(C_OUTPUT_FIFO_66_DMWIDTH),
        .C_OUTPUT_FIFO_67_DMWIDTH(C_OUTPUT_FIFO_67_DMWIDTH),
        .C_OUTPUT_FIFO_68_DMWIDTH(C_OUTPUT_FIFO_68_DMWIDTH),
        .C_OUTPUT_FIFO_69_DMWIDTH(C_OUTPUT_FIFO_69_DMWIDTH),
        .C_OUTPUT_FIFO_70_DMWIDTH(C_OUTPUT_FIFO_70_DMWIDTH),
        .C_OUTPUT_FIFO_71_DMWIDTH(C_OUTPUT_FIFO_71_DMWIDTH),
        .C_OUTPUT_FIFO_72_DMWIDTH(C_OUTPUT_FIFO_72_DMWIDTH),
        .C_OUTPUT_FIFO_73_DMWIDTH(C_OUTPUT_FIFO_73_DMWIDTH),
        .C_OUTPUT_FIFO_74_DMWIDTH(C_OUTPUT_FIFO_74_DMWIDTH),
        .C_OUTPUT_FIFO_75_DMWIDTH(C_OUTPUT_FIFO_75_DMWIDTH),
        .C_OUTPUT_FIFO_76_DMWIDTH(C_OUTPUT_FIFO_76_DMWIDTH),
        .C_OUTPUT_FIFO_77_DMWIDTH(C_OUTPUT_FIFO_77_DMWIDTH),
        .C_OUTPUT_FIFO_78_DMWIDTH(C_OUTPUT_FIFO_78_DMWIDTH),
        .C_OUTPUT_FIFO_79_DMWIDTH(C_OUTPUT_FIFO_79_DMWIDTH),
        .C_OUTPUT_FIFO_80_DMWIDTH(C_OUTPUT_FIFO_80_DMWIDTH),
        .C_OUTPUT_FIFO_81_DMWIDTH(C_OUTPUT_FIFO_81_DMWIDTH),
        .C_OUTPUT_FIFO_82_DMWIDTH(C_OUTPUT_FIFO_82_DMWIDTH),
        .C_OUTPUT_FIFO_83_DMWIDTH(C_OUTPUT_FIFO_83_DMWIDTH),
        .C_OUTPUT_FIFO_84_DMWIDTH(C_OUTPUT_FIFO_84_DMWIDTH),
        .C_OUTPUT_FIFO_85_DMWIDTH(C_OUTPUT_FIFO_85_DMWIDTH),
        .C_OUTPUT_FIFO_86_DMWIDTH(C_OUTPUT_FIFO_86_DMWIDTH),
        .C_OUTPUT_FIFO_87_DMWIDTH(C_OUTPUT_FIFO_87_DMWIDTH),
        .C_OUTPUT_FIFO_88_DMWIDTH(C_OUTPUT_FIFO_88_DMWIDTH),
        .C_OUTPUT_FIFO_89_DMWIDTH(C_OUTPUT_FIFO_89_DMWIDTH),
        .C_OUTPUT_FIFO_90_DMWIDTH(C_OUTPUT_FIFO_90_DMWIDTH),
        .C_OUTPUT_FIFO_91_DMWIDTH(C_OUTPUT_FIFO_91_DMWIDTH),
        .C_OUTPUT_FIFO_92_DMWIDTH(C_OUTPUT_FIFO_92_DMWIDTH),
        .C_OUTPUT_FIFO_93_DMWIDTH(C_OUTPUT_FIFO_93_DMWIDTH),
        .C_OUTPUT_FIFO_94_DMWIDTH(C_OUTPUT_FIFO_94_DMWIDTH),
        .C_OUTPUT_FIFO_95_DMWIDTH(C_OUTPUT_FIFO_95_DMWIDTH),
        .C_OUTPUT_FIFO_96_DMWIDTH(C_OUTPUT_FIFO_96_DMWIDTH),
        .C_OUTPUT_FIFO_97_DMWIDTH(C_OUTPUT_FIFO_97_DMWIDTH),
        .C_OUTPUT_FIFO_98_DMWIDTH(C_OUTPUT_FIFO_98_DMWIDTH),
        .C_OUTPUT_FIFO_99_DMWIDTH(C_OUTPUT_FIFO_99_DMWIDTH),
        .C_OUTPUT_FIFO_100_DMWIDTH(C_OUTPUT_FIFO_100_DMWIDTH),
        .C_OUTPUT_FIFO_101_DMWIDTH(C_OUTPUT_FIFO_101_DMWIDTH),
        .C_OUTPUT_FIFO_102_DMWIDTH(C_OUTPUT_FIFO_102_DMWIDTH),
        .C_OUTPUT_FIFO_103_DMWIDTH(C_OUTPUT_FIFO_103_DMWIDTH),
        .C_OUTPUT_FIFO_104_DMWIDTH(C_OUTPUT_FIFO_104_DMWIDTH),
        .C_OUTPUT_FIFO_105_DMWIDTH(C_OUTPUT_FIFO_105_DMWIDTH),
        .C_OUTPUT_FIFO_106_DMWIDTH(C_OUTPUT_FIFO_106_DMWIDTH),
        .C_OUTPUT_FIFO_107_DMWIDTH(C_OUTPUT_FIFO_107_DMWIDTH),
        .C_OUTPUT_FIFO_108_DMWIDTH(C_OUTPUT_FIFO_108_DMWIDTH),
        .C_OUTPUT_FIFO_109_DMWIDTH(C_OUTPUT_FIFO_109_DMWIDTH),
        .C_OUTPUT_FIFO_110_DMWIDTH(C_OUTPUT_FIFO_110_DMWIDTH),
        .C_OUTPUT_FIFO_111_DMWIDTH(C_OUTPUT_FIFO_111_DMWIDTH),
        .C_OUTPUT_FIFO_112_DMWIDTH(C_OUTPUT_FIFO_112_DMWIDTH),
        .C_OUTPUT_FIFO_113_DMWIDTH(C_OUTPUT_FIFO_113_DMWIDTH),
        .C_OUTPUT_FIFO_114_DMWIDTH(C_OUTPUT_FIFO_114_DMWIDTH),
        .C_OUTPUT_FIFO_115_DMWIDTH(C_OUTPUT_FIFO_115_DMWIDTH),
        .C_OUTPUT_FIFO_116_DMWIDTH(C_OUTPUT_FIFO_116_DMWIDTH),
        .C_OUTPUT_FIFO_117_DMWIDTH(C_OUTPUT_FIFO_117_DMWIDTH),
        .C_OUTPUT_FIFO_118_DMWIDTH(C_OUTPUT_FIFO_118_DMWIDTH),
        .C_OUTPUT_FIFO_119_DMWIDTH(C_OUTPUT_FIFO_119_DMWIDTH),
        .C_OUTPUT_FIFO_120_DMWIDTH(C_OUTPUT_FIFO_120_DMWIDTH),
        .C_OUTPUT_FIFO_121_DMWIDTH(C_OUTPUT_FIFO_121_DMWIDTH),
        .C_OUTPUT_FIFO_122_DMWIDTH(C_OUTPUT_FIFO_122_DMWIDTH),
        .C_OUTPUT_FIFO_123_DMWIDTH(C_OUTPUT_FIFO_123_DMWIDTH),
        .C_OUTPUT_FIFO_124_DMWIDTH(C_OUTPUT_FIFO_124_DMWIDTH),
        .C_OUTPUT_FIFO_125_DMWIDTH(C_OUTPUT_FIFO_125_DMWIDTH),
        .C_OUTPUT_FIFO_126_DMWIDTH(C_OUTPUT_FIFO_126_DMWIDTH),
        .C_OUTPUT_FIFO_127_DMWIDTH(C_OUTPUT_FIFO_127_DMWIDTH)
    ) out_fifo_args_i (
        .acc_clk(aclk),
        .dm_clk(s_axi_aclk),
        .aresetn(s_axi_aresetn),
        .out_fifo_allow(outfifo_ctrl_allow),
        .m_axis_fifo_0_tlast(m_axis_fifo_0_tlast),
        .m_axis_fifo_0_tvalid(m_axis_fifo_0_tvalid),
        .m_axis_fifo_0_tkeep(m_axis_fifo_0_tkeep),
        .m_axis_fifo_0_tstrb(m_axis_fifo_0_tstrb),
        .m_axis_fifo_0_tdata(m_axis_fifo_0_tdata),
        .m_axis_fifo_0_tready(m_axis_fifo_0_tready),
        .ap_fifo_oarg_0_full_n(ap_fifo_oarg_0_full_n),
        .ap_fifo_oarg_0_din(ap_fifo_oarg_0_din),
        .ap_fifo_oarg_0_write(ap_fifo_oarg_0_write),
        .m_axis_fifo_1_tlast(m_axis_fifo_1_tlast),
        .m_axis_fifo_1_tvalid(m_axis_fifo_1_tvalid),
        .m_axis_fifo_1_tkeep(m_axis_fifo_1_tkeep),
        .m_axis_fifo_1_tstrb(m_axis_fifo_1_tstrb),
        .m_axis_fifo_1_tdata(m_axis_fifo_1_tdata),
        .m_axis_fifo_1_tready(m_axis_fifo_1_tready),
        .ap_fifo_oarg_1_full_n(ap_fifo_oarg_1_full_n),
        .ap_fifo_oarg_1_din(ap_fifo_oarg_1_din),
        .ap_fifo_oarg_1_write(ap_fifo_oarg_1_write),
        .m_axis_fifo_2_tlast(m_axis_fifo_2_tlast),
        .m_axis_fifo_2_tvalid(m_axis_fifo_2_tvalid),
        .m_axis_fifo_2_tkeep(m_axis_fifo_2_tkeep),
        .m_axis_fifo_2_tstrb(m_axis_fifo_2_tstrb),
        .m_axis_fifo_2_tdata(m_axis_fifo_2_tdata),
        .m_axis_fifo_2_tready(m_axis_fifo_2_tready),
        .ap_fifo_oarg_2_full_n(ap_fifo_oarg_2_full_n),
        .ap_fifo_oarg_2_din(ap_fifo_oarg_2_din),
        .ap_fifo_oarg_2_write(ap_fifo_oarg_2_write),
        .m_axis_fifo_3_tlast(m_axis_fifo_3_tlast),
        .m_axis_fifo_3_tvalid(m_axis_fifo_3_tvalid),
        .m_axis_fifo_3_tkeep(m_axis_fifo_3_tkeep),
        .m_axis_fifo_3_tstrb(m_axis_fifo_3_tstrb),
        .m_axis_fifo_3_tdata(m_axis_fifo_3_tdata),
        .m_axis_fifo_3_tready(m_axis_fifo_3_tready),
        .ap_fifo_oarg_3_full_n(ap_fifo_oarg_3_full_n),
        .ap_fifo_oarg_3_din(ap_fifo_oarg_3_din),
        .ap_fifo_oarg_3_write(ap_fifo_oarg_3_write),
        .m_axis_fifo_4_tlast(m_axis_fifo_4_tlast),
        .m_axis_fifo_4_tvalid(m_axis_fifo_4_tvalid),
        .m_axis_fifo_4_tkeep(m_axis_fifo_4_tkeep),
        .m_axis_fifo_4_tstrb(m_axis_fifo_4_tstrb),
        .m_axis_fifo_4_tdata(m_axis_fifo_4_tdata),
        .m_axis_fifo_4_tready(m_axis_fifo_4_tready),
        .ap_fifo_oarg_4_full_n(ap_fifo_oarg_4_full_n),
        .ap_fifo_oarg_4_din(ap_fifo_oarg_4_din),
        .ap_fifo_oarg_4_write(ap_fifo_oarg_4_write),
        .m_axis_fifo_5_tlast(m_axis_fifo_5_tlast),
        .m_axis_fifo_5_tvalid(m_axis_fifo_5_tvalid),
        .m_axis_fifo_5_tkeep(m_axis_fifo_5_tkeep),
        .m_axis_fifo_5_tstrb(m_axis_fifo_5_tstrb),
        .m_axis_fifo_5_tdata(m_axis_fifo_5_tdata),
        .m_axis_fifo_5_tready(m_axis_fifo_5_tready),
        .ap_fifo_oarg_5_full_n(ap_fifo_oarg_5_full_n),
        .ap_fifo_oarg_5_din(ap_fifo_oarg_5_din),
        .ap_fifo_oarg_5_write(ap_fifo_oarg_5_write),
        .m_axis_fifo_6_tlast(m_axis_fifo_6_tlast),
        .m_axis_fifo_6_tvalid(m_axis_fifo_6_tvalid),
        .m_axis_fifo_6_tkeep(m_axis_fifo_6_tkeep),
        .m_axis_fifo_6_tstrb(m_axis_fifo_6_tstrb),
        .m_axis_fifo_6_tdata(m_axis_fifo_6_tdata),
        .m_axis_fifo_6_tready(m_axis_fifo_6_tready),
        .ap_fifo_oarg_6_full_n(ap_fifo_oarg_6_full_n),
        .ap_fifo_oarg_6_din(ap_fifo_oarg_6_din),
        .ap_fifo_oarg_6_write(ap_fifo_oarg_6_write),
        .m_axis_fifo_7_tlast(m_axis_fifo_7_tlast),
        .m_axis_fifo_7_tvalid(m_axis_fifo_7_tvalid),
        .m_axis_fifo_7_tkeep(m_axis_fifo_7_tkeep),
        .m_axis_fifo_7_tstrb(m_axis_fifo_7_tstrb),
        .m_axis_fifo_7_tdata(m_axis_fifo_7_tdata),
        .m_axis_fifo_7_tready(m_axis_fifo_7_tready),
        .ap_fifo_oarg_7_full_n(ap_fifo_oarg_7_full_n),
        .ap_fifo_oarg_7_din(ap_fifo_oarg_7_din),
        .ap_fifo_oarg_7_write(ap_fifo_oarg_7_write),
        .m_axis_fifo_8_tlast(m_axis_fifo_8_tlast),
        .m_axis_fifo_8_tvalid(m_axis_fifo_8_tvalid),
        .m_axis_fifo_8_tkeep(m_axis_fifo_8_tkeep),
        .m_axis_fifo_8_tstrb(m_axis_fifo_8_tstrb),
        .m_axis_fifo_8_tdata(m_axis_fifo_8_tdata),
        .m_axis_fifo_8_tready(m_axis_fifo_8_tready),
        .ap_fifo_oarg_8_full_n(ap_fifo_oarg_8_full_n),
        .ap_fifo_oarg_8_din(ap_fifo_oarg_8_din),
        .ap_fifo_oarg_8_write(ap_fifo_oarg_8_write),
        .m_axis_fifo_9_tlast(m_axis_fifo_9_tlast),
        .m_axis_fifo_9_tvalid(m_axis_fifo_9_tvalid),
        .m_axis_fifo_9_tkeep(m_axis_fifo_9_tkeep),
        .m_axis_fifo_9_tstrb(m_axis_fifo_9_tstrb),
        .m_axis_fifo_9_tdata(m_axis_fifo_9_tdata),
        .m_axis_fifo_9_tready(m_axis_fifo_9_tready),
        .ap_fifo_oarg_9_full_n(ap_fifo_oarg_9_full_n),
        .ap_fifo_oarg_9_din(ap_fifo_oarg_9_din),
        .ap_fifo_oarg_9_write(ap_fifo_oarg_9_write),
        .m_axis_fifo_10_tlast(m_axis_fifo_10_tlast),
        .m_axis_fifo_10_tvalid(m_axis_fifo_10_tvalid),
        .m_axis_fifo_10_tkeep(m_axis_fifo_10_tkeep),
        .m_axis_fifo_10_tstrb(m_axis_fifo_10_tstrb),
        .m_axis_fifo_10_tdata(m_axis_fifo_10_tdata),
        .m_axis_fifo_10_tready(m_axis_fifo_10_tready),
        .ap_fifo_oarg_10_full_n(ap_fifo_oarg_10_full_n),
        .ap_fifo_oarg_10_din(ap_fifo_oarg_10_din),
        .ap_fifo_oarg_10_write(ap_fifo_oarg_10_write),
        .m_axis_fifo_11_tlast(m_axis_fifo_11_tlast),
        .m_axis_fifo_11_tvalid(m_axis_fifo_11_tvalid),
        .m_axis_fifo_11_tkeep(m_axis_fifo_11_tkeep),
        .m_axis_fifo_11_tstrb(m_axis_fifo_11_tstrb),
        .m_axis_fifo_11_tdata(m_axis_fifo_11_tdata),
        .m_axis_fifo_11_tready(m_axis_fifo_11_tready),
        .ap_fifo_oarg_11_full_n(ap_fifo_oarg_11_full_n),
        .ap_fifo_oarg_11_din(ap_fifo_oarg_11_din),
        .ap_fifo_oarg_11_write(ap_fifo_oarg_11_write),
        .m_axis_fifo_12_tlast(m_axis_fifo_12_tlast),
        .m_axis_fifo_12_tvalid(m_axis_fifo_12_tvalid),
        .m_axis_fifo_12_tkeep(m_axis_fifo_12_tkeep),
        .m_axis_fifo_12_tstrb(m_axis_fifo_12_tstrb),
        .m_axis_fifo_12_tdata(m_axis_fifo_12_tdata),
        .m_axis_fifo_12_tready(m_axis_fifo_12_tready),
        .ap_fifo_oarg_12_full_n(ap_fifo_oarg_12_full_n),
        .ap_fifo_oarg_12_din(ap_fifo_oarg_12_din),
        .ap_fifo_oarg_12_write(ap_fifo_oarg_12_write),
        .m_axis_fifo_13_tlast(m_axis_fifo_13_tlast),
        .m_axis_fifo_13_tvalid(m_axis_fifo_13_tvalid),
        .m_axis_fifo_13_tkeep(m_axis_fifo_13_tkeep),
        .m_axis_fifo_13_tstrb(m_axis_fifo_13_tstrb),
        .m_axis_fifo_13_tdata(m_axis_fifo_13_tdata),
        .m_axis_fifo_13_tready(m_axis_fifo_13_tready),
        .ap_fifo_oarg_13_full_n(ap_fifo_oarg_13_full_n),
        .ap_fifo_oarg_13_din(ap_fifo_oarg_13_din),
        .ap_fifo_oarg_13_write(ap_fifo_oarg_13_write),
        .m_axis_fifo_14_tlast(m_axis_fifo_14_tlast),
        .m_axis_fifo_14_tvalid(m_axis_fifo_14_tvalid),
        .m_axis_fifo_14_tkeep(m_axis_fifo_14_tkeep),
        .m_axis_fifo_14_tstrb(m_axis_fifo_14_tstrb),
        .m_axis_fifo_14_tdata(m_axis_fifo_14_tdata),
        .m_axis_fifo_14_tready(m_axis_fifo_14_tready),
        .ap_fifo_oarg_14_full_n(ap_fifo_oarg_14_full_n),
        .ap_fifo_oarg_14_din(ap_fifo_oarg_14_din),
        .ap_fifo_oarg_14_write(ap_fifo_oarg_14_write),
        .m_axis_fifo_15_tlast(m_axis_fifo_15_tlast),
        .m_axis_fifo_15_tvalid(m_axis_fifo_15_tvalid),
        .m_axis_fifo_15_tkeep(m_axis_fifo_15_tkeep),
        .m_axis_fifo_15_tstrb(m_axis_fifo_15_tstrb),
        .m_axis_fifo_15_tdata(m_axis_fifo_15_tdata),
        .m_axis_fifo_15_tready(m_axis_fifo_15_tready),
        .ap_fifo_oarg_15_full_n(ap_fifo_oarg_15_full_n),
        .ap_fifo_oarg_15_din(ap_fifo_oarg_15_din),
        .ap_fifo_oarg_15_write(ap_fifo_oarg_15_write),
        .m_axis_fifo_16_tlast(m_axis_fifo_16_tlast),
        .m_axis_fifo_16_tvalid(m_axis_fifo_16_tvalid),
        .m_axis_fifo_16_tkeep(m_axis_fifo_16_tkeep),
        .m_axis_fifo_16_tstrb(m_axis_fifo_16_tstrb),
        .m_axis_fifo_16_tdata(m_axis_fifo_16_tdata),
        .m_axis_fifo_16_tready(m_axis_fifo_16_tready),
        .ap_fifo_oarg_16_full_n(ap_fifo_oarg_16_full_n),
        .ap_fifo_oarg_16_din(ap_fifo_oarg_16_din),
        .ap_fifo_oarg_16_write(ap_fifo_oarg_16_write),
        .m_axis_fifo_17_tlast(m_axis_fifo_17_tlast),
        .m_axis_fifo_17_tvalid(m_axis_fifo_17_tvalid),
        .m_axis_fifo_17_tkeep(m_axis_fifo_17_tkeep),
        .m_axis_fifo_17_tstrb(m_axis_fifo_17_tstrb),
        .m_axis_fifo_17_tdata(m_axis_fifo_17_tdata),
        .m_axis_fifo_17_tready(m_axis_fifo_17_tready),
        .ap_fifo_oarg_17_full_n(ap_fifo_oarg_17_full_n),
        .ap_fifo_oarg_17_din(ap_fifo_oarg_17_din),
        .ap_fifo_oarg_17_write(ap_fifo_oarg_17_write),
        .m_axis_fifo_18_tlast(m_axis_fifo_18_tlast),
        .m_axis_fifo_18_tvalid(m_axis_fifo_18_tvalid),
        .m_axis_fifo_18_tkeep(m_axis_fifo_18_tkeep),
        .m_axis_fifo_18_tstrb(m_axis_fifo_18_tstrb),
        .m_axis_fifo_18_tdata(m_axis_fifo_18_tdata),
        .m_axis_fifo_18_tready(m_axis_fifo_18_tready),
        .ap_fifo_oarg_18_full_n(ap_fifo_oarg_18_full_n),
        .ap_fifo_oarg_18_din(ap_fifo_oarg_18_din),
        .ap_fifo_oarg_18_write(ap_fifo_oarg_18_write),
        .m_axis_fifo_19_tlast(m_axis_fifo_19_tlast),
        .m_axis_fifo_19_tvalid(m_axis_fifo_19_tvalid),
        .m_axis_fifo_19_tkeep(m_axis_fifo_19_tkeep),
        .m_axis_fifo_19_tstrb(m_axis_fifo_19_tstrb),
        .m_axis_fifo_19_tdata(m_axis_fifo_19_tdata),
        .m_axis_fifo_19_tready(m_axis_fifo_19_tready),
        .ap_fifo_oarg_19_full_n(ap_fifo_oarg_19_full_n),
        .ap_fifo_oarg_19_din(ap_fifo_oarg_19_din),
        .ap_fifo_oarg_19_write(ap_fifo_oarg_19_write),
        .m_axis_fifo_20_tlast(m_axis_fifo_20_tlast),
        .m_axis_fifo_20_tvalid(m_axis_fifo_20_tvalid),
        .m_axis_fifo_20_tkeep(m_axis_fifo_20_tkeep),
        .m_axis_fifo_20_tstrb(m_axis_fifo_20_tstrb),
        .m_axis_fifo_20_tdata(m_axis_fifo_20_tdata),
        .m_axis_fifo_20_tready(m_axis_fifo_20_tready),
        .ap_fifo_oarg_20_full_n(ap_fifo_oarg_20_full_n),
        .ap_fifo_oarg_20_din(ap_fifo_oarg_20_din),
        .ap_fifo_oarg_20_write(ap_fifo_oarg_20_write),
        .m_axis_fifo_21_tlast(m_axis_fifo_21_tlast),
        .m_axis_fifo_21_tvalid(m_axis_fifo_21_tvalid),
        .m_axis_fifo_21_tkeep(m_axis_fifo_21_tkeep),
        .m_axis_fifo_21_tstrb(m_axis_fifo_21_tstrb),
        .m_axis_fifo_21_tdata(m_axis_fifo_21_tdata),
        .m_axis_fifo_21_tready(m_axis_fifo_21_tready),
        .ap_fifo_oarg_21_full_n(ap_fifo_oarg_21_full_n),
        .ap_fifo_oarg_21_din(ap_fifo_oarg_21_din),
        .ap_fifo_oarg_21_write(ap_fifo_oarg_21_write),
        .m_axis_fifo_22_tlast(m_axis_fifo_22_tlast),
        .m_axis_fifo_22_tvalid(m_axis_fifo_22_tvalid),
        .m_axis_fifo_22_tkeep(m_axis_fifo_22_tkeep),
        .m_axis_fifo_22_tstrb(m_axis_fifo_22_tstrb),
        .m_axis_fifo_22_tdata(m_axis_fifo_22_tdata),
        .m_axis_fifo_22_tready(m_axis_fifo_22_tready),
        .ap_fifo_oarg_22_full_n(ap_fifo_oarg_22_full_n),
        .ap_fifo_oarg_22_din(ap_fifo_oarg_22_din),
        .ap_fifo_oarg_22_write(ap_fifo_oarg_22_write),
        .m_axis_fifo_23_tlast(m_axis_fifo_23_tlast),
        .m_axis_fifo_23_tvalid(m_axis_fifo_23_tvalid),
        .m_axis_fifo_23_tkeep(m_axis_fifo_23_tkeep),
        .m_axis_fifo_23_tstrb(m_axis_fifo_23_tstrb),
        .m_axis_fifo_23_tdata(m_axis_fifo_23_tdata),
        .m_axis_fifo_23_tready(m_axis_fifo_23_tready),
        .ap_fifo_oarg_23_full_n(ap_fifo_oarg_23_full_n),
        .ap_fifo_oarg_23_din(ap_fifo_oarg_23_din),
        .ap_fifo_oarg_23_write(ap_fifo_oarg_23_write),
        .m_axis_fifo_24_tlast(m_axis_fifo_24_tlast),
        .m_axis_fifo_24_tvalid(m_axis_fifo_24_tvalid),
        .m_axis_fifo_24_tkeep(m_axis_fifo_24_tkeep),
        .m_axis_fifo_24_tstrb(m_axis_fifo_24_tstrb),
        .m_axis_fifo_24_tdata(m_axis_fifo_24_tdata),
        .m_axis_fifo_24_tready(m_axis_fifo_24_tready),
        .ap_fifo_oarg_24_full_n(ap_fifo_oarg_24_full_n),
        .ap_fifo_oarg_24_din(ap_fifo_oarg_24_din),
        .ap_fifo_oarg_24_write(ap_fifo_oarg_24_write),
        .m_axis_fifo_25_tlast(m_axis_fifo_25_tlast),
        .m_axis_fifo_25_tvalid(m_axis_fifo_25_tvalid),
        .m_axis_fifo_25_tkeep(m_axis_fifo_25_tkeep),
        .m_axis_fifo_25_tstrb(m_axis_fifo_25_tstrb),
        .m_axis_fifo_25_tdata(m_axis_fifo_25_tdata),
        .m_axis_fifo_25_tready(m_axis_fifo_25_tready),
        .ap_fifo_oarg_25_full_n(ap_fifo_oarg_25_full_n),
        .ap_fifo_oarg_25_din(ap_fifo_oarg_25_din),
        .ap_fifo_oarg_25_write(ap_fifo_oarg_25_write),
        .m_axis_fifo_26_tlast(m_axis_fifo_26_tlast),
        .m_axis_fifo_26_tvalid(m_axis_fifo_26_tvalid),
        .m_axis_fifo_26_tkeep(m_axis_fifo_26_tkeep),
        .m_axis_fifo_26_tstrb(m_axis_fifo_26_tstrb),
        .m_axis_fifo_26_tdata(m_axis_fifo_26_tdata),
        .m_axis_fifo_26_tready(m_axis_fifo_26_tready),
        .ap_fifo_oarg_26_full_n(ap_fifo_oarg_26_full_n),
        .ap_fifo_oarg_26_din(ap_fifo_oarg_26_din),
        .ap_fifo_oarg_26_write(ap_fifo_oarg_26_write),
        .m_axis_fifo_27_tlast(m_axis_fifo_27_tlast),
        .m_axis_fifo_27_tvalid(m_axis_fifo_27_tvalid),
        .m_axis_fifo_27_tkeep(m_axis_fifo_27_tkeep),
        .m_axis_fifo_27_tstrb(m_axis_fifo_27_tstrb),
        .m_axis_fifo_27_tdata(m_axis_fifo_27_tdata),
        .m_axis_fifo_27_tready(m_axis_fifo_27_tready),
        .ap_fifo_oarg_27_full_n(ap_fifo_oarg_27_full_n),
        .ap_fifo_oarg_27_din(ap_fifo_oarg_27_din),
        .ap_fifo_oarg_27_write(ap_fifo_oarg_27_write),
        .m_axis_fifo_28_tlast(m_axis_fifo_28_tlast),
        .m_axis_fifo_28_tvalid(m_axis_fifo_28_tvalid),
        .m_axis_fifo_28_tkeep(m_axis_fifo_28_tkeep),
        .m_axis_fifo_28_tstrb(m_axis_fifo_28_tstrb),
        .m_axis_fifo_28_tdata(m_axis_fifo_28_tdata),
        .m_axis_fifo_28_tready(m_axis_fifo_28_tready),
        .ap_fifo_oarg_28_full_n(ap_fifo_oarg_28_full_n),
        .ap_fifo_oarg_28_din(ap_fifo_oarg_28_din),
        .ap_fifo_oarg_28_write(ap_fifo_oarg_28_write),
        .m_axis_fifo_29_tlast(m_axis_fifo_29_tlast),
        .m_axis_fifo_29_tvalid(m_axis_fifo_29_tvalid),
        .m_axis_fifo_29_tkeep(m_axis_fifo_29_tkeep),
        .m_axis_fifo_29_tstrb(m_axis_fifo_29_tstrb),
        .m_axis_fifo_29_tdata(m_axis_fifo_29_tdata),
        .m_axis_fifo_29_tready(m_axis_fifo_29_tready),
        .ap_fifo_oarg_29_full_n(ap_fifo_oarg_29_full_n),
        .ap_fifo_oarg_29_din(ap_fifo_oarg_29_din),
        .ap_fifo_oarg_29_write(ap_fifo_oarg_29_write),
        .m_axis_fifo_30_tlast(m_axis_fifo_30_tlast),
        .m_axis_fifo_30_tvalid(m_axis_fifo_30_tvalid),
        .m_axis_fifo_30_tkeep(m_axis_fifo_30_tkeep),
        .m_axis_fifo_30_tstrb(m_axis_fifo_30_tstrb),
        .m_axis_fifo_30_tdata(m_axis_fifo_30_tdata),
        .m_axis_fifo_30_tready(m_axis_fifo_30_tready),
        .ap_fifo_oarg_30_full_n(ap_fifo_oarg_30_full_n),
        .ap_fifo_oarg_30_din(ap_fifo_oarg_30_din),
        .ap_fifo_oarg_30_write(ap_fifo_oarg_30_write),
        .m_axis_fifo_31_tlast(m_axis_fifo_31_tlast),
        .m_axis_fifo_31_tvalid(m_axis_fifo_31_tvalid),
        .m_axis_fifo_31_tkeep(m_axis_fifo_31_tkeep),
        .m_axis_fifo_31_tstrb(m_axis_fifo_31_tstrb),
        .m_axis_fifo_31_tdata(m_axis_fifo_31_tdata),
        .m_axis_fifo_31_tready(m_axis_fifo_31_tready),
        .ap_fifo_oarg_31_full_n(ap_fifo_oarg_31_full_n),
        .ap_fifo_oarg_31_din(ap_fifo_oarg_31_din),
        .ap_fifo_oarg_31_write(ap_fifo_oarg_31_write),
        .m_axis_fifo_32_tlast(m_axis_fifo_32_tlast),
        .m_axis_fifo_32_tvalid(m_axis_fifo_32_tvalid),
        .m_axis_fifo_32_tkeep(m_axis_fifo_32_tkeep),
        .m_axis_fifo_32_tstrb(m_axis_fifo_32_tstrb),
        .m_axis_fifo_32_tdata(m_axis_fifo_32_tdata),
        .m_axis_fifo_32_tready(m_axis_fifo_32_tready),
        .ap_fifo_oarg_32_full_n(ap_fifo_oarg_32_full_n),
        .ap_fifo_oarg_32_din(ap_fifo_oarg_32_din),
        .ap_fifo_oarg_32_write(ap_fifo_oarg_32_write),
        .m_axis_fifo_33_tlast(m_axis_fifo_33_tlast),
        .m_axis_fifo_33_tvalid(m_axis_fifo_33_tvalid),
        .m_axis_fifo_33_tkeep(m_axis_fifo_33_tkeep),
        .m_axis_fifo_33_tstrb(m_axis_fifo_33_tstrb),
        .m_axis_fifo_33_tdata(m_axis_fifo_33_tdata),
        .m_axis_fifo_33_tready(m_axis_fifo_33_tready),
        .ap_fifo_oarg_33_full_n(ap_fifo_oarg_33_full_n),
        .ap_fifo_oarg_33_din(ap_fifo_oarg_33_din),
        .ap_fifo_oarg_33_write(ap_fifo_oarg_33_write),
        .m_axis_fifo_34_tlast(m_axis_fifo_34_tlast),
        .m_axis_fifo_34_tvalid(m_axis_fifo_34_tvalid),
        .m_axis_fifo_34_tkeep(m_axis_fifo_34_tkeep),
        .m_axis_fifo_34_tstrb(m_axis_fifo_34_tstrb),
        .m_axis_fifo_34_tdata(m_axis_fifo_34_tdata),
        .m_axis_fifo_34_tready(m_axis_fifo_34_tready),
        .ap_fifo_oarg_34_full_n(ap_fifo_oarg_34_full_n),
        .ap_fifo_oarg_34_din(ap_fifo_oarg_34_din),
        .ap_fifo_oarg_34_write(ap_fifo_oarg_34_write),
        .m_axis_fifo_35_tlast(m_axis_fifo_35_tlast),
        .m_axis_fifo_35_tvalid(m_axis_fifo_35_tvalid),
        .m_axis_fifo_35_tkeep(m_axis_fifo_35_tkeep),
        .m_axis_fifo_35_tstrb(m_axis_fifo_35_tstrb),
        .m_axis_fifo_35_tdata(m_axis_fifo_35_tdata),
        .m_axis_fifo_35_tready(m_axis_fifo_35_tready),
        .ap_fifo_oarg_35_full_n(ap_fifo_oarg_35_full_n),
        .ap_fifo_oarg_35_din(ap_fifo_oarg_35_din),
        .ap_fifo_oarg_35_write(ap_fifo_oarg_35_write),
        .m_axis_fifo_36_tlast(m_axis_fifo_36_tlast),
        .m_axis_fifo_36_tvalid(m_axis_fifo_36_tvalid),
        .m_axis_fifo_36_tkeep(m_axis_fifo_36_tkeep),
        .m_axis_fifo_36_tstrb(m_axis_fifo_36_tstrb),
        .m_axis_fifo_36_tdata(m_axis_fifo_36_tdata),
        .m_axis_fifo_36_tready(m_axis_fifo_36_tready),
        .ap_fifo_oarg_36_full_n(ap_fifo_oarg_36_full_n),
        .ap_fifo_oarg_36_din(ap_fifo_oarg_36_din),
        .ap_fifo_oarg_36_write(ap_fifo_oarg_36_write),
        .m_axis_fifo_37_tlast(m_axis_fifo_37_tlast),
        .m_axis_fifo_37_tvalid(m_axis_fifo_37_tvalid),
        .m_axis_fifo_37_tkeep(m_axis_fifo_37_tkeep),
        .m_axis_fifo_37_tstrb(m_axis_fifo_37_tstrb),
        .m_axis_fifo_37_tdata(m_axis_fifo_37_tdata),
        .m_axis_fifo_37_tready(m_axis_fifo_37_tready),
        .ap_fifo_oarg_37_full_n(ap_fifo_oarg_37_full_n),
        .ap_fifo_oarg_37_din(ap_fifo_oarg_37_din),
        .ap_fifo_oarg_37_write(ap_fifo_oarg_37_write),
        .m_axis_fifo_38_tlast(m_axis_fifo_38_tlast),
        .m_axis_fifo_38_tvalid(m_axis_fifo_38_tvalid),
        .m_axis_fifo_38_tkeep(m_axis_fifo_38_tkeep),
        .m_axis_fifo_38_tstrb(m_axis_fifo_38_tstrb),
        .m_axis_fifo_38_tdata(m_axis_fifo_38_tdata),
        .m_axis_fifo_38_tready(m_axis_fifo_38_tready),
        .ap_fifo_oarg_38_full_n(ap_fifo_oarg_38_full_n),
        .ap_fifo_oarg_38_din(ap_fifo_oarg_38_din),
        .ap_fifo_oarg_38_write(ap_fifo_oarg_38_write),
        .m_axis_fifo_39_tlast(m_axis_fifo_39_tlast),
        .m_axis_fifo_39_tvalid(m_axis_fifo_39_tvalid),
        .m_axis_fifo_39_tkeep(m_axis_fifo_39_tkeep),
        .m_axis_fifo_39_tstrb(m_axis_fifo_39_tstrb),
        .m_axis_fifo_39_tdata(m_axis_fifo_39_tdata),
        .m_axis_fifo_39_tready(m_axis_fifo_39_tready),
        .ap_fifo_oarg_39_full_n(ap_fifo_oarg_39_full_n),
        .ap_fifo_oarg_39_din(ap_fifo_oarg_39_din),
        .ap_fifo_oarg_39_write(ap_fifo_oarg_39_write),
        .m_axis_fifo_40_tlast(m_axis_fifo_40_tlast),
        .m_axis_fifo_40_tvalid(m_axis_fifo_40_tvalid),
        .m_axis_fifo_40_tkeep(m_axis_fifo_40_tkeep),
        .m_axis_fifo_40_tstrb(m_axis_fifo_40_tstrb),
        .m_axis_fifo_40_tdata(m_axis_fifo_40_tdata),
        .m_axis_fifo_40_tready(m_axis_fifo_40_tready),
        .ap_fifo_oarg_40_full_n(ap_fifo_oarg_40_full_n),
        .ap_fifo_oarg_40_din(ap_fifo_oarg_40_din),
        .ap_fifo_oarg_40_write(ap_fifo_oarg_40_write),
        .m_axis_fifo_41_tlast(m_axis_fifo_41_tlast),
        .m_axis_fifo_41_tvalid(m_axis_fifo_41_tvalid),
        .m_axis_fifo_41_tkeep(m_axis_fifo_41_tkeep),
        .m_axis_fifo_41_tstrb(m_axis_fifo_41_tstrb),
        .m_axis_fifo_41_tdata(m_axis_fifo_41_tdata),
        .m_axis_fifo_41_tready(m_axis_fifo_41_tready),
        .ap_fifo_oarg_41_full_n(ap_fifo_oarg_41_full_n),
        .ap_fifo_oarg_41_din(ap_fifo_oarg_41_din),
        .ap_fifo_oarg_41_write(ap_fifo_oarg_41_write),
        .m_axis_fifo_42_tlast(m_axis_fifo_42_tlast),
        .m_axis_fifo_42_tvalid(m_axis_fifo_42_tvalid),
        .m_axis_fifo_42_tkeep(m_axis_fifo_42_tkeep),
        .m_axis_fifo_42_tstrb(m_axis_fifo_42_tstrb),
        .m_axis_fifo_42_tdata(m_axis_fifo_42_tdata),
        .m_axis_fifo_42_tready(m_axis_fifo_42_tready),
        .ap_fifo_oarg_42_full_n(ap_fifo_oarg_42_full_n),
        .ap_fifo_oarg_42_din(ap_fifo_oarg_42_din),
        .ap_fifo_oarg_42_write(ap_fifo_oarg_42_write),
        .m_axis_fifo_43_tlast(m_axis_fifo_43_tlast),
        .m_axis_fifo_43_tvalid(m_axis_fifo_43_tvalid),
        .m_axis_fifo_43_tkeep(m_axis_fifo_43_tkeep),
        .m_axis_fifo_43_tstrb(m_axis_fifo_43_tstrb),
        .m_axis_fifo_43_tdata(m_axis_fifo_43_tdata),
        .m_axis_fifo_43_tready(m_axis_fifo_43_tready),
        .ap_fifo_oarg_43_full_n(ap_fifo_oarg_43_full_n),
        .ap_fifo_oarg_43_din(ap_fifo_oarg_43_din),
        .ap_fifo_oarg_43_write(ap_fifo_oarg_43_write),
        .m_axis_fifo_44_tlast(m_axis_fifo_44_tlast),
        .m_axis_fifo_44_tvalid(m_axis_fifo_44_tvalid),
        .m_axis_fifo_44_tkeep(m_axis_fifo_44_tkeep),
        .m_axis_fifo_44_tstrb(m_axis_fifo_44_tstrb),
        .m_axis_fifo_44_tdata(m_axis_fifo_44_tdata),
        .m_axis_fifo_44_tready(m_axis_fifo_44_tready),
        .ap_fifo_oarg_44_full_n(ap_fifo_oarg_44_full_n),
        .ap_fifo_oarg_44_din(ap_fifo_oarg_44_din),
        .ap_fifo_oarg_44_write(ap_fifo_oarg_44_write),
        .m_axis_fifo_45_tlast(m_axis_fifo_45_tlast),
        .m_axis_fifo_45_tvalid(m_axis_fifo_45_tvalid),
        .m_axis_fifo_45_tkeep(m_axis_fifo_45_tkeep),
        .m_axis_fifo_45_tstrb(m_axis_fifo_45_tstrb),
        .m_axis_fifo_45_tdata(m_axis_fifo_45_tdata),
        .m_axis_fifo_45_tready(m_axis_fifo_45_tready),
        .ap_fifo_oarg_45_full_n(ap_fifo_oarg_45_full_n),
        .ap_fifo_oarg_45_din(ap_fifo_oarg_45_din),
        .ap_fifo_oarg_45_write(ap_fifo_oarg_45_write),
        .m_axis_fifo_46_tlast(m_axis_fifo_46_tlast),
        .m_axis_fifo_46_tvalid(m_axis_fifo_46_tvalid),
        .m_axis_fifo_46_tkeep(m_axis_fifo_46_tkeep),
        .m_axis_fifo_46_tstrb(m_axis_fifo_46_tstrb),
        .m_axis_fifo_46_tdata(m_axis_fifo_46_tdata),
        .m_axis_fifo_46_tready(m_axis_fifo_46_tready),
        .ap_fifo_oarg_46_full_n(ap_fifo_oarg_46_full_n),
        .ap_fifo_oarg_46_din(ap_fifo_oarg_46_din),
        .ap_fifo_oarg_46_write(ap_fifo_oarg_46_write),
        .m_axis_fifo_47_tlast(m_axis_fifo_47_tlast),
        .m_axis_fifo_47_tvalid(m_axis_fifo_47_tvalid),
        .m_axis_fifo_47_tkeep(m_axis_fifo_47_tkeep),
        .m_axis_fifo_47_tstrb(m_axis_fifo_47_tstrb),
        .m_axis_fifo_47_tdata(m_axis_fifo_47_tdata),
        .m_axis_fifo_47_tready(m_axis_fifo_47_tready),
        .ap_fifo_oarg_47_full_n(ap_fifo_oarg_47_full_n),
        .ap_fifo_oarg_47_din(ap_fifo_oarg_47_din),
        .ap_fifo_oarg_47_write(ap_fifo_oarg_47_write),
        .m_axis_fifo_48_tlast(m_axis_fifo_48_tlast),
        .m_axis_fifo_48_tvalid(m_axis_fifo_48_tvalid),
        .m_axis_fifo_48_tkeep(m_axis_fifo_48_tkeep),
        .m_axis_fifo_48_tstrb(m_axis_fifo_48_tstrb),
        .m_axis_fifo_48_tdata(m_axis_fifo_48_tdata),
        .m_axis_fifo_48_tready(m_axis_fifo_48_tready),
        .ap_fifo_oarg_48_full_n(ap_fifo_oarg_48_full_n),
        .ap_fifo_oarg_48_din(ap_fifo_oarg_48_din),
        .ap_fifo_oarg_48_write(ap_fifo_oarg_48_write),
        .m_axis_fifo_49_tlast(m_axis_fifo_49_tlast),
        .m_axis_fifo_49_tvalid(m_axis_fifo_49_tvalid),
        .m_axis_fifo_49_tkeep(m_axis_fifo_49_tkeep),
        .m_axis_fifo_49_tstrb(m_axis_fifo_49_tstrb),
        .m_axis_fifo_49_tdata(m_axis_fifo_49_tdata),
        .m_axis_fifo_49_tready(m_axis_fifo_49_tready),
        .ap_fifo_oarg_49_full_n(ap_fifo_oarg_49_full_n),
        .ap_fifo_oarg_49_din(ap_fifo_oarg_49_din),
        .ap_fifo_oarg_49_write(ap_fifo_oarg_49_write),
        .m_axis_fifo_50_tlast(m_axis_fifo_50_tlast),
        .m_axis_fifo_50_tvalid(m_axis_fifo_50_tvalid),
        .m_axis_fifo_50_tkeep(m_axis_fifo_50_tkeep),
        .m_axis_fifo_50_tstrb(m_axis_fifo_50_tstrb),
        .m_axis_fifo_50_tdata(m_axis_fifo_50_tdata),
        .m_axis_fifo_50_tready(m_axis_fifo_50_tready),
        .ap_fifo_oarg_50_full_n(ap_fifo_oarg_50_full_n),
        .ap_fifo_oarg_50_din(ap_fifo_oarg_50_din),
        .ap_fifo_oarg_50_write(ap_fifo_oarg_50_write),
        .m_axis_fifo_51_tlast(m_axis_fifo_51_tlast),
        .m_axis_fifo_51_tvalid(m_axis_fifo_51_tvalid),
        .m_axis_fifo_51_tkeep(m_axis_fifo_51_tkeep),
        .m_axis_fifo_51_tstrb(m_axis_fifo_51_tstrb),
        .m_axis_fifo_51_tdata(m_axis_fifo_51_tdata),
        .m_axis_fifo_51_tready(m_axis_fifo_51_tready),
        .ap_fifo_oarg_51_full_n(ap_fifo_oarg_51_full_n),
        .ap_fifo_oarg_51_din(ap_fifo_oarg_51_din),
        .ap_fifo_oarg_51_write(ap_fifo_oarg_51_write),
        .m_axis_fifo_52_tlast(m_axis_fifo_52_tlast),
        .m_axis_fifo_52_tvalid(m_axis_fifo_52_tvalid),
        .m_axis_fifo_52_tkeep(m_axis_fifo_52_tkeep),
        .m_axis_fifo_52_tstrb(m_axis_fifo_52_tstrb),
        .m_axis_fifo_52_tdata(m_axis_fifo_52_tdata),
        .m_axis_fifo_52_tready(m_axis_fifo_52_tready),
        .ap_fifo_oarg_52_full_n(ap_fifo_oarg_52_full_n),
        .ap_fifo_oarg_52_din(ap_fifo_oarg_52_din),
        .ap_fifo_oarg_52_write(ap_fifo_oarg_52_write),
        .m_axis_fifo_53_tlast(m_axis_fifo_53_tlast),
        .m_axis_fifo_53_tvalid(m_axis_fifo_53_tvalid),
        .m_axis_fifo_53_tkeep(m_axis_fifo_53_tkeep),
        .m_axis_fifo_53_tstrb(m_axis_fifo_53_tstrb),
        .m_axis_fifo_53_tdata(m_axis_fifo_53_tdata),
        .m_axis_fifo_53_tready(m_axis_fifo_53_tready),
        .ap_fifo_oarg_53_full_n(ap_fifo_oarg_53_full_n),
        .ap_fifo_oarg_53_din(ap_fifo_oarg_53_din),
        .ap_fifo_oarg_53_write(ap_fifo_oarg_53_write),
        .m_axis_fifo_54_tlast(m_axis_fifo_54_tlast),
        .m_axis_fifo_54_tvalid(m_axis_fifo_54_tvalid),
        .m_axis_fifo_54_tkeep(m_axis_fifo_54_tkeep),
        .m_axis_fifo_54_tstrb(m_axis_fifo_54_tstrb),
        .m_axis_fifo_54_tdata(m_axis_fifo_54_tdata),
        .m_axis_fifo_54_tready(m_axis_fifo_54_tready),
        .ap_fifo_oarg_54_full_n(ap_fifo_oarg_54_full_n),
        .ap_fifo_oarg_54_din(ap_fifo_oarg_54_din),
        .ap_fifo_oarg_54_write(ap_fifo_oarg_54_write),
        .m_axis_fifo_55_tlast(m_axis_fifo_55_tlast),
        .m_axis_fifo_55_tvalid(m_axis_fifo_55_tvalid),
        .m_axis_fifo_55_tkeep(m_axis_fifo_55_tkeep),
        .m_axis_fifo_55_tstrb(m_axis_fifo_55_tstrb),
        .m_axis_fifo_55_tdata(m_axis_fifo_55_tdata),
        .m_axis_fifo_55_tready(m_axis_fifo_55_tready),
        .ap_fifo_oarg_55_full_n(ap_fifo_oarg_55_full_n),
        .ap_fifo_oarg_55_din(ap_fifo_oarg_55_din),
        .ap_fifo_oarg_55_write(ap_fifo_oarg_55_write),
        .m_axis_fifo_56_tlast(m_axis_fifo_56_tlast),
        .m_axis_fifo_56_tvalid(m_axis_fifo_56_tvalid),
        .m_axis_fifo_56_tkeep(m_axis_fifo_56_tkeep),
        .m_axis_fifo_56_tstrb(m_axis_fifo_56_tstrb),
        .m_axis_fifo_56_tdata(m_axis_fifo_56_tdata),
        .m_axis_fifo_56_tready(m_axis_fifo_56_tready),
        .ap_fifo_oarg_56_full_n(ap_fifo_oarg_56_full_n),
        .ap_fifo_oarg_56_din(ap_fifo_oarg_56_din),
        .ap_fifo_oarg_56_write(ap_fifo_oarg_56_write),
        .m_axis_fifo_57_tlast(m_axis_fifo_57_tlast),
        .m_axis_fifo_57_tvalid(m_axis_fifo_57_tvalid),
        .m_axis_fifo_57_tkeep(m_axis_fifo_57_tkeep),
        .m_axis_fifo_57_tstrb(m_axis_fifo_57_tstrb),
        .m_axis_fifo_57_tdata(m_axis_fifo_57_tdata),
        .m_axis_fifo_57_tready(m_axis_fifo_57_tready),
        .ap_fifo_oarg_57_full_n(ap_fifo_oarg_57_full_n),
        .ap_fifo_oarg_57_din(ap_fifo_oarg_57_din),
        .ap_fifo_oarg_57_write(ap_fifo_oarg_57_write),
        .m_axis_fifo_58_tlast(m_axis_fifo_58_tlast),
        .m_axis_fifo_58_tvalid(m_axis_fifo_58_tvalid),
        .m_axis_fifo_58_tkeep(m_axis_fifo_58_tkeep),
        .m_axis_fifo_58_tstrb(m_axis_fifo_58_tstrb),
        .m_axis_fifo_58_tdata(m_axis_fifo_58_tdata),
        .m_axis_fifo_58_tready(m_axis_fifo_58_tready),
        .ap_fifo_oarg_58_full_n(ap_fifo_oarg_58_full_n),
        .ap_fifo_oarg_58_din(ap_fifo_oarg_58_din),
        .ap_fifo_oarg_58_write(ap_fifo_oarg_58_write),
        .m_axis_fifo_59_tlast(m_axis_fifo_59_tlast),
        .m_axis_fifo_59_tvalid(m_axis_fifo_59_tvalid),
        .m_axis_fifo_59_tkeep(m_axis_fifo_59_tkeep),
        .m_axis_fifo_59_tstrb(m_axis_fifo_59_tstrb),
        .m_axis_fifo_59_tdata(m_axis_fifo_59_tdata),
        .m_axis_fifo_59_tready(m_axis_fifo_59_tready),
        .ap_fifo_oarg_59_full_n(ap_fifo_oarg_59_full_n),
        .ap_fifo_oarg_59_din(ap_fifo_oarg_59_din),
        .ap_fifo_oarg_59_write(ap_fifo_oarg_59_write),
        .m_axis_fifo_60_tlast(m_axis_fifo_60_tlast),
        .m_axis_fifo_60_tvalid(m_axis_fifo_60_tvalid),
        .m_axis_fifo_60_tkeep(m_axis_fifo_60_tkeep),
        .m_axis_fifo_60_tstrb(m_axis_fifo_60_tstrb),
        .m_axis_fifo_60_tdata(m_axis_fifo_60_tdata),
        .m_axis_fifo_60_tready(m_axis_fifo_60_tready),
        .ap_fifo_oarg_60_full_n(ap_fifo_oarg_60_full_n),
        .ap_fifo_oarg_60_din(ap_fifo_oarg_60_din),
        .ap_fifo_oarg_60_write(ap_fifo_oarg_60_write),
        .m_axis_fifo_61_tlast(m_axis_fifo_61_tlast),
        .m_axis_fifo_61_tvalid(m_axis_fifo_61_tvalid),
        .m_axis_fifo_61_tkeep(m_axis_fifo_61_tkeep),
        .m_axis_fifo_61_tstrb(m_axis_fifo_61_tstrb),
        .m_axis_fifo_61_tdata(m_axis_fifo_61_tdata),
        .m_axis_fifo_61_tready(m_axis_fifo_61_tready),
        .ap_fifo_oarg_61_full_n(ap_fifo_oarg_61_full_n),
        .ap_fifo_oarg_61_din(ap_fifo_oarg_61_din),
        .ap_fifo_oarg_61_write(ap_fifo_oarg_61_write),
        .m_axis_fifo_62_tlast(m_axis_fifo_62_tlast),
        .m_axis_fifo_62_tvalid(m_axis_fifo_62_tvalid),
        .m_axis_fifo_62_tkeep(m_axis_fifo_62_tkeep),
        .m_axis_fifo_62_tstrb(m_axis_fifo_62_tstrb),
        .m_axis_fifo_62_tdata(m_axis_fifo_62_tdata),
        .m_axis_fifo_62_tready(m_axis_fifo_62_tready),
        .ap_fifo_oarg_62_full_n(ap_fifo_oarg_62_full_n),
        .ap_fifo_oarg_62_din(ap_fifo_oarg_62_din),
        .ap_fifo_oarg_62_write(ap_fifo_oarg_62_write),
        .m_axis_fifo_63_tlast(m_axis_fifo_63_tlast),
        .m_axis_fifo_63_tvalid(m_axis_fifo_63_tvalid),
        .m_axis_fifo_63_tkeep(m_axis_fifo_63_tkeep),
        .m_axis_fifo_63_tstrb(m_axis_fifo_63_tstrb),
        .m_axis_fifo_63_tdata(m_axis_fifo_63_tdata),
        .m_axis_fifo_63_tready(m_axis_fifo_63_tready),
        .ap_fifo_oarg_63_full_n(ap_fifo_oarg_63_full_n),
        .ap_fifo_oarg_63_din(ap_fifo_oarg_63_din),
        .ap_fifo_oarg_63_write(ap_fifo_oarg_63_write),
        .m_axis_fifo_64_tlast(m_axis_fifo_64_tlast),
        .m_axis_fifo_64_tvalid(m_axis_fifo_64_tvalid),
        .m_axis_fifo_64_tkeep(m_axis_fifo_64_tkeep),
        .m_axis_fifo_64_tstrb(m_axis_fifo_64_tstrb),
        .m_axis_fifo_64_tdata(m_axis_fifo_64_tdata),
        .m_axis_fifo_64_tready(m_axis_fifo_64_tready),
        .ap_fifo_oarg_64_full_n(ap_fifo_oarg_64_full_n),
        .ap_fifo_oarg_64_din(ap_fifo_oarg_64_din),
        .ap_fifo_oarg_64_write(ap_fifo_oarg_64_write),
        .m_axis_fifo_65_tlast(m_axis_fifo_65_tlast),
        .m_axis_fifo_65_tvalid(m_axis_fifo_65_tvalid),
        .m_axis_fifo_65_tkeep(m_axis_fifo_65_tkeep),
        .m_axis_fifo_65_tstrb(m_axis_fifo_65_tstrb),
        .m_axis_fifo_65_tdata(m_axis_fifo_65_tdata),
        .m_axis_fifo_65_tready(m_axis_fifo_65_tready),
        .ap_fifo_oarg_65_full_n(ap_fifo_oarg_65_full_n),
        .ap_fifo_oarg_65_din(ap_fifo_oarg_65_din),
        .ap_fifo_oarg_65_write(ap_fifo_oarg_65_write),
        .m_axis_fifo_66_tlast(m_axis_fifo_66_tlast),
        .m_axis_fifo_66_tvalid(m_axis_fifo_66_tvalid),
        .m_axis_fifo_66_tkeep(m_axis_fifo_66_tkeep),
        .m_axis_fifo_66_tstrb(m_axis_fifo_66_tstrb),
        .m_axis_fifo_66_tdata(m_axis_fifo_66_tdata),
        .m_axis_fifo_66_tready(m_axis_fifo_66_tready),
        .ap_fifo_oarg_66_full_n(ap_fifo_oarg_66_full_n),
        .ap_fifo_oarg_66_din(ap_fifo_oarg_66_din),
        .ap_fifo_oarg_66_write(ap_fifo_oarg_66_write),
        .m_axis_fifo_67_tlast(m_axis_fifo_67_tlast),
        .m_axis_fifo_67_tvalid(m_axis_fifo_67_tvalid),
        .m_axis_fifo_67_tkeep(m_axis_fifo_67_tkeep),
        .m_axis_fifo_67_tstrb(m_axis_fifo_67_tstrb),
        .m_axis_fifo_67_tdata(m_axis_fifo_67_tdata),
        .m_axis_fifo_67_tready(m_axis_fifo_67_tready),
        .ap_fifo_oarg_67_full_n(ap_fifo_oarg_67_full_n),
        .ap_fifo_oarg_67_din(ap_fifo_oarg_67_din),
        .ap_fifo_oarg_67_write(ap_fifo_oarg_67_write),
        .m_axis_fifo_68_tlast(m_axis_fifo_68_tlast),
        .m_axis_fifo_68_tvalid(m_axis_fifo_68_tvalid),
        .m_axis_fifo_68_tkeep(m_axis_fifo_68_tkeep),
        .m_axis_fifo_68_tstrb(m_axis_fifo_68_tstrb),
        .m_axis_fifo_68_tdata(m_axis_fifo_68_tdata),
        .m_axis_fifo_68_tready(m_axis_fifo_68_tready),
        .ap_fifo_oarg_68_full_n(ap_fifo_oarg_68_full_n),
        .ap_fifo_oarg_68_din(ap_fifo_oarg_68_din),
        .ap_fifo_oarg_68_write(ap_fifo_oarg_68_write),
        .m_axis_fifo_69_tlast(m_axis_fifo_69_tlast),
        .m_axis_fifo_69_tvalid(m_axis_fifo_69_tvalid),
        .m_axis_fifo_69_tkeep(m_axis_fifo_69_tkeep),
        .m_axis_fifo_69_tstrb(m_axis_fifo_69_tstrb),
        .m_axis_fifo_69_tdata(m_axis_fifo_69_tdata),
        .m_axis_fifo_69_tready(m_axis_fifo_69_tready),
        .ap_fifo_oarg_69_full_n(ap_fifo_oarg_69_full_n),
        .ap_fifo_oarg_69_din(ap_fifo_oarg_69_din),
        .ap_fifo_oarg_69_write(ap_fifo_oarg_69_write),
        .m_axis_fifo_70_tlast(m_axis_fifo_70_tlast),
        .m_axis_fifo_70_tvalid(m_axis_fifo_70_tvalid),
        .m_axis_fifo_70_tkeep(m_axis_fifo_70_tkeep),
        .m_axis_fifo_70_tstrb(m_axis_fifo_70_tstrb),
        .m_axis_fifo_70_tdata(m_axis_fifo_70_tdata),
        .m_axis_fifo_70_tready(m_axis_fifo_70_tready),
        .ap_fifo_oarg_70_full_n(ap_fifo_oarg_70_full_n),
        .ap_fifo_oarg_70_din(ap_fifo_oarg_70_din),
        .ap_fifo_oarg_70_write(ap_fifo_oarg_70_write),
        .m_axis_fifo_71_tlast(m_axis_fifo_71_tlast),
        .m_axis_fifo_71_tvalid(m_axis_fifo_71_tvalid),
        .m_axis_fifo_71_tkeep(m_axis_fifo_71_tkeep),
        .m_axis_fifo_71_tstrb(m_axis_fifo_71_tstrb),
        .m_axis_fifo_71_tdata(m_axis_fifo_71_tdata),
        .m_axis_fifo_71_tready(m_axis_fifo_71_tready),
        .ap_fifo_oarg_71_full_n(ap_fifo_oarg_71_full_n),
        .ap_fifo_oarg_71_din(ap_fifo_oarg_71_din),
        .ap_fifo_oarg_71_write(ap_fifo_oarg_71_write),
        .m_axis_fifo_72_tlast(m_axis_fifo_72_tlast),
        .m_axis_fifo_72_tvalid(m_axis_fifo_72_tvalid),
        .m_axis_fifo_72_tkeep(m_axis_fifo_72_tkeep),
        .m_axis_fifo_72_tstrb(m_axis_fifo_72_tstrb),
        .m_axis_fifo_72_tdata(m_axis_fifo_72_tdata),
        .m_axis_fifo_72_tready(m_axis_fifo_72_tready),
        .ap_fifo_oarg_72_full_n(ap_fifo_oarg_72_full_n),
        .ap_fifo_oarg_72_din(ap_fifo_oarg_72_din),
        .ap_fifo_oarg_72_write(ap_fifo_oarg_72_write),
        .m_axis_fifo_73_tlast(m_axis_fifo_73_tlast),
        .m_axis_fifo_73_tvalid(m_axis_fifo_73_tvalid),
        .m_axis_fifo_73_tkeep(m_axis_fifo_73_tkeep),
        .m_axis_fifo_73_tstrb(m_axis_fifo_73_tstrb),
        .m_axis_fifo_73_tdata(m_axis_fifo_73_tdata),
        .m_axis_fifo_73_tready(m_axis_fifo_73_tready),
        .ap_fifo_oarg_73_full_n(ap_fifo_oarg_73_full_n),
        .ap_fifo_oarg_73_din(ap_fifo_oarg_73_din),
        .ap_fifo_oarg_73_write(ap_fifo_oarg_73_write),
        .m_axis_fifo_74_tlast(m_axis_fifo_74_tlast),
        .m_axis_fifo_74_tvalid(m_axis_fifo_74_tvalid),
        .m_axis_fifo_74_tkeep(m_axis_fifo_74_tkeep),
        .m_axis_fifo_74_tstrb(m_axis_fifo_74_tstrb),
        .m_axis_fifo_74_tdata(m_axis_fifo_74_tdata),
        .m_axis_fifo_74_tready(m_axis_fifo_74_tready),
        .ap_fifo_oarg_74_full_n(ap_fifo_oarg_74_full_n),
        .ap_fifo_oarg_74_din(ap_fifo_oarg_74_din),
        .ap_fifo_oarg_74_write(ap_fifo_oarg_74_write),
        .m_axis_fifo_75_tlast(m_axis_fifo_75_tlast),
        .m_axis_fifo_75_tvalid(m_axis_fifo_75_tvalid),
        .m_axis_fifo_75_tkeep(m_axis_fifo_75_tkeep),
        .m_axis_fifo_75_tstrb(m_axis_fifo_75_tstrb),
        .m_axis_fifo_75_tdata(m_axis_fifo_75_tdata),
        .m_axis_fifo_75_tready(m_axis_fifo_75_tready),
        .ap_fifo_oarg_75_full_n(ap_fifo_oarg_75_full_n),
        .ap_fifo_oarg_75_din(ap_fifo_oarg_75_din),
        .ap_fifo_oarg_75_write(ap_fifo_oarg_75_write),
        .m_axis_fifo_76_tlast(m_axis_fifo_76_tlast),
        .m_axis_fifo_76_tvalid(m_axis_fifo_76_tvalid),
        .m_axis_fifo_76_tkeep(m_axis_fifo_76_tkeep),
        .m_axis_fifo_76_tstrb(m_axis_fifo_76_tstrb),
        .m_axis_fifo_76_tdata(m_axis_fifo_76_tdata),
        .m_axis_fifo_76_tready(m_axis_fifo_76_tready),
        .ap_fifo_oarg_76_full_n(ap_fifo_oarg_76_full_n),
        .ap_fifo_oarg_76_din(ap_fifo_oarg_76_din),
        .ap_fifo_oarg_76_write(ap_fifo_oarg_76_write),
        .m_axis_fifo_77_tlast(m_axis_fifo_77_tlast),
        .m_axis_fifo_77_tvalid(m_axis_fifo_77_tvalid),
        .m_axis_fifo_77_tkeep(m_axis_fifo_77_tkeep),
        .m_axis_fifo_77_tstrb(m_axis_fifo_77_tstrb),
        .m_axis_fifo_77_tdata(m_axis_fifo_77_tdata),
        .m_axis_fifo_77_tready(m_axis_fifo_77_tready),
        .ap_fifo_oarg_77_full_n(ap_fifo_oarg_77_full_n),
        .ap_fifo_oarg_77_din(ap_fifo_oarg_77_din),
        .ap_fifo_oarg_77_write(ap_fifo_oarg_77_write),
        .m_axis_fifo_78_tlast(m_axis_fifo_78_tlast),
        .m_axis_fifo_78_tvalid(m_axis_fifo_78_tvalid),
        .m_axis_fifo_78_tkeep(m_axis_fifo_78_tkeep),
        .m_axis_fifo_78_tstrb(m_axis_fifo_78_tstrb),
        .m_axis_fifo_78_tdata(m_axis_fifo_78_tdata),
        .m_axis_fifo_78_tready(m_axis_fifo_78_tready),
        .ap_fifo_oarg_78_full_n(ap_fifo_oarg_78_full_n),
        .ap_fifo_oarg_78_din(ap_fifo_oarg_78_din),
        .ap_fifo_oarg_78_write(ap_fifo_oarg_78_write),
        .m_axis_fifo_79_tlast(m_axis_fifo_79_tlast),
        .m_axis_fifo_79_tvalid(m_axis_fifo_79_tvalid),
        .m_axis_fifo_79_tkeep(m_axis_fifo_79_tkeep),
        .m_axis_fifo_79_tstrb(m_axis_fifo_79_tstrb),
        .m_axis_fifo_79_tdata(m_axis_fifo_79_tdata),
        .m_axis_fifo_79_tready(m_axis_fifo_79_tready),
        .ap_fifo_oarg_79_full_n(ap_fifo_oarg_79_full_n),
        .ap_fifo_oarg_79_din(ap_fifo_oarg_79_din),
        .ap_fifo_oarg_79_write(ap_fifo_oarg_79_write),
        .m_axis_fifo_80_tlast(m_axis_fifo_80_tlast),
        .m_axis_fifo_80_tvalid(m_axis_fifo_80_tvalid),
        .m_axis_fifo_80_tkeep(m_axis_fifo_80_tkeep),
        .m_axis_fifo_80_tstrb(m_axis_fifo_80_tstrb),
        .m_axis_fifo_80_tdata(m_axis_fifo_80_tdata),
        .m_axis_fifo_80_tready(m_axis_fifo_80_tready),
        .ap_fifo_oarg_80_full_n(ap_fifo_oarg_80_full_n),
        .ap_fifo_oarg_80_din(ap_fifo_oarg_80_din),
        .ap_fifo_oarg_80_write(ap_fifo_oarg_80_write),
        .m_axis_fifo_81_tlast(m_axis_fifo_81_tlast),
        .m_axis_fifo_81_tvalid(m_axis_fifo_81_tvalid),
        .m_axis_fifo_81_tkeep(m_axis_fifo_81_tkeep),
        .m_axis_fifo_81_tstrb(m_axis_fifo_81_tstrb),
        .m_axis_fifo_81_tdata(m_axis_fifo_81_tdata),
        .m_axis_fifo_81_tready(m_axis_fifo_81_tready),
        .ap_fifo_oarg_81_full_n(ap_fifo_oarg_81_full_n),
        .ap_fifo_oarg_81_din(ap_fifo_oarg_81_din),
        .ap_fifo_oarg_81_write(ap_fifo_oarg_81_write),
        .m_axis_fifo_82_tlast(m_axis_fifo_82_tlast),
        .m_axis_fifo_82_tvalid(m_axis_fifo_82_tvalid),
        .m_axis_fifo_82_tkeep(m_axis_fifo_82_tkeep),
        .m_axis_fifo_82_tstrb(m_axis_fifo_82_tstrb),
        .m_axis_fifo_82_tdata(m_axis_fifo_82_tdata),
        .m_axis_fifo_82_tready(m_axis_fifo_82_tready),
        .ap_fifo_oarg_82_full_n(ap_fifo_oarg_82_full_n),
        .ap_fifo_oarg_82_din(ap_fifo_oarg_82_din),
        .ap_fifo_oarg_82_write(ap_fifo_oarg_82_write),
        .m_axis_fifo_83_tlast(m_axis_fifo_83_tlast),
        .m_axis_fifo_83_tvalid(m_axis_fifo_83_tvalid),
        .m_axis_fifo_83_tkeep(m_axis_fifo_83_tkeep),
        .m_axis_fifo_83_tstrb(m_axis_fifo_83_tstrb),
        .m_axis_fifo_83_tdata(m_axis_fifo_83_tdata),
        .m_axis_fifo_83_tready(m_axis_fifo_83_tready),
        .ap_fifo_oarg_83_full_n(ap_fifo_oarg_83_full_n),
        .ap_fifo_oarg_83_din(ap_fifo_oarg_83_din),
        .ap_fifo_oarg_83_write(ap_fifo_oarg_83_write),
        .m_axis_fifo_84_tlast(m_axis_fifo_84_tlast),
        .m_axis_fifo_84_tvalid(m_axis_fifo_84_tvalid),
        .m_axis_fifo_84_tkeep(m_axis_fifo_84_tkeep),
        .m_axis_fifo_84_tstrb(m_axis_fifo_84_tstrb),
        .m_axis_fifo_84_tdata(m_axis_fifo_84_tdata),
        .m_axis_fifo_84_tready(m_axis_fifo_84_tready),
        .ap_fifo_oarg_84_full_n(ap_fifo_oarg_84_full_n),
        .ap_fifo_oarg_84_din(ap_fifo_oarg_84_din),
        .ap_fifo_oarg_84_write(ap_fifo_oarg_84_write),
        .m_axis_fifo_85_tlast(m_axis_fifo_85_tlast),
        .m_axis_fifo_85_tvalid(m_axis_fifo_85_tvalid),
        .m_axis_fifo_85_tkeep(m_axis_fifo_85_tkeep),
        .m_axis_fifo_85_tstrb(m_axis_fifo_85_tstrb),
        .m_axis_fifo_85_tdata(m_axis_fifo_85_tdata),
        .m_axis_fifo_85_tready(m_axis_fifo_85_tready),
        .ap_fifo_oarg_85_full_n(ap_fifo_oarg_85_full_n),
        .ap_fifo_oarg_85_din(ap_fifo_oarg_85_din),
        .ap_fifo_oarg_85_write(ap_fifo_oarg_85_write),
        .m_axis_fifo_86_tlast(m_axis_fifo_86_tlast),
        .m_axis_fifo_86_tvalid(m_axis_fifo_86_tvalid),
        .m_axis_fifo_86_tkeep(m_axis_fifo_86_tkeep),
        .m_axis_fifo_86_tstrb(m_axis_fifo_86_tstrb),
        .m_axis_fifo_86_tdata(m_axis_fifo_86_tdata),
        .m_axis_fifo_86_tready(m_axis_fifo_86_tready),
        .ap_fifo_oarg_86_full_n(ap_fifo_oarg_86_full_n),
        .ap_fifo_oarg_86_din(ap_fifo_oarg_86_din),
        .ap_fifo_oarg_86_write(ap_fifo_oarg_86_write),
        .m_axis_fifo_87_tlast(m_axis_fifo_87_tlast),
        .m_axis_fifo_87_tvalid(m_axis_fifo_87_tvalid),
        .m_axis_fifo_87_tkeep(m_axis_fifo_87_tkeep),
        .m_axis_fifo_87_tstrb(m_axis_fifo_87_tstrb),
        .m_axis_fifo_87_tdata(m_axis_fifo_87_tdata),
        .m_axis_fifo_87_tready(m_axis_fifo_87_tready),
        .ap_fifo_oarg_87_full_n(ap_fifo_oarg_87_full_n),
        .ap_fifo_oarg_87_din(ap_fifo_oarg_87_din),
        .ap_fifo_oarg_87_write(ap_fifo_oarg_87_write),
        .m_axis_fifo_88_tlast(m_axis_fifo_88_tlast),
        .m_axis_fifo_88_tvalid(m_axis_fifo_88_tvalid),
        .m_axis_fifo_88_tkeep(m_axis_fifo_88_tkeep),
        .m_axis_fifo_88_tstrb(m_axis_fifo_88_tstrb),
        .m_axis_fifo_88_tdata(m_axis_fifo_88_tdata),
        .m_axis_fifo_88_tready(m_axis_fifo_88_tready),
        .ap_fifo_oarg_88_full_n(ap_fifo_oarg_88_full_n),
        .ap_fifo_oarg_88_din(ap_fifo_oarg_88_din),
        .ap_fifo_oarg_88_write(ap_fifo_oarg_88_write),
        .m_axis_fifo_89_tlast(m_axis_fifo_89_tlast),
        .m_axis_fifo_89_tvalid(m_axis_fifo_89_tvalid),
        .m_axis_fifo_89_tkeep(m_axis_fifo_89_tkeep),
        .m_axis_fifo_89_tstrb(m_axis_fifo_89_tstrb),
        .m_axis_fifo_89_tdata(m_axis_fifo_89_tdata),
        .m_axis_fifo_89_tready(m_axis_fifo_89_tready),
        .ap_fifo_oarg_89_full_n(ap_fifo_oarg_89_full_n),
        .ap_fifo_oarg_89_din(ap_fifo_oarg_89_din),
        .ap_fifo_oarg_89_write(ap_fifo_oarg_89_write),
        .m_axis_fifo_90_tlast(m_axis_fifo_90_tlast),
        .m_axis_fifo_90_tvalid(m_axis_fifo_90_tvalid),
        .m_axis_fifo_90_tkeep(m_axis_fifo_90_tkeep),
        .m_axis_fifo_90_tstrb(m_axis_fifo_90_tstrb),
        .m_axis_fifo_90_tdata(m_axis_fifo_90_tdata),
        .m_axis_fifo_90_tready(m_axis_fifo_90_tready),
        .ap_fifo_oarg_90_full_n(ap_fifo_oarg_90_full_n),
        .ap_fifo_oarg_90_din(ap_fifo_oarg_90_din),
        .ap_fifo_oarg_90_write(ap_fifo_oarg_90_write),
        .m_axis_fifo_91_tlast(m_axis_fifo_91_tlast),
        .m_axis_fifo_91_tvalid(m_axis_fifo_91_tvalid),
        .m_axis_fifo_91_tkeep(m_axis_fifo_91_tkeep),
        .m_axis_fifo_91_tstrb(m_axis_fifo_91_tstrb),
        .m_axis_fifo_91_tdata(m_axis_fifo_91_tdata),
        .m_axis_fifo_91_tready(m_axis_fifo_91_tready),
        .ap_fifo_oarg_91_full_n(ap_fifo_oarg_91_full_n),
        .ap_fifo_oarg_91_din(ap_fifo_oarg_91_din),
        .ap_fifo_oarg_91_write(ap_fifo_oarg_91_write),
        .m_axis_fifo_92_tlast(m_axis_fifo_92_tlast),
        .m_axis_fifo_92_tvalid(m_axis_fifo_92_tvalid),
        .m_axis_fifo_92_tkeep(m_axis_fifo_92_tkeep),
        .m_axis_fifo_92_tstrb(m_axis_fifo_92_tstrb),
        .m_axis_fifo_92_tdata(m_axis_fifo_92_tdata),
        .m_axis_fifo_92_tready(m_axis_fifo_92_tready),
        .ap_fifo_oarg_92_full_n(ap_fifo_oarg_92_full_n),
        .ap_fifo_oarg_92_din(ap_fifo_oarg_92_din),
        .ap_fifo_oarg_92_write(ap_fifo_oarg_92_write),
        .m_axis_fifo_93_tlast(m_axis_fifo_93_tlast),
        .m_axis_fifo_93_tvalid(m_axis_fifo_93_tvalid),
        .m_axis_fifo_93_tkeep(m_axis_fifo_93_tkeep),
        .m_axis_fifo_93_tstrb(m_axis_fifo_93_tstrb),
        .m_axis_fifo_93_tdata(m_axis_fifo_93_tdata),
        .m_axis_fifo_93_tready(m_axis_fifo_93_tready),
        .ap_fifo_oarg_93_full_n(ap_fifo_oarg_93_full_n),
        .ap_fifo_oarg_93_din(ap_fifo_oarg_93_din),
        .ap_fifo_oarg_93_write(ap_fifo_oarg_93_write),
        .m_axis_fifo_94_tlast(m_axis_fifo_94_tlast),
        .m_axis_fifo_94_tvalid(m_axis_fifo_94_tvalid),
        .m_axis_fifo_94_tkeep(m_axis_fifo_94_tkeep),
        .m_axis_fifo_94_tstrb(m_axis_fifo_94_tstrb),
        .m_axis_fifo_94_tdata(m_axis_fifo_94_tdata),
        .m_axis_fifo_94_tready(m_axis_fifo_94_tready),
        .ap_fifo_oarg_94_full_n(ap_fifo_oarg_94_full_n),
        .ap_fifo_oarg_94_din(ap_fifo_oarg_94_din),
        .ap_fifo_oarg_94_write(ap_fifo_oarg_94_write),
        .m_axis_fifo_95_tlast(m_axis_fifo_95_tlast),
        .m_axis_fifo_95_tvalid(m_axis_fifo_95_tvalid),
        .m_axis_fifo_95_tkeep(m_axis_fifo_95_tkeep),
        .m_axis_fifo_95_tstrb(m_axis_fifo_95_tstrb),
        .m_axis_fifo_95_tdata(m_axis_fifo_95_tdata),
        .m_axis_fifo_95_tready(m_axis_fifo_95_tready),
        .ap_fifo_oarg_95_full_n(ap_fifo_oarg_95_full_n),
        .ap_fifo_oarg_95_din(ap_fifo_oarg_95_din),
        .ap_fifo_oarg_95_write(ap_fifo_oarg_95_write),
        .m_axis_fifo_96_tlast(m_axis_fifo_96_tlast),
        .m_axis_fifo_96_tvalid(m_axis_fifo_96_tvalid),
        .m_axis_fifo_96_tkeep(m_axis_fifo_96_tkeep),
        .m_axis_fifo_96_tstrb(m_axis_fifo_96_tstrb),
        .m_axis_fifo_96_tdata(m_axis_fifo_96_tdata),
        .m_axis_fifo_96_tready(m_axis_fifo_96_tready),
        .ap_fifo_oarg_96_full_n(ap_fifo_oarg_96_full_n),
        .ap_fifo_oarg_96_din(ap_fifo_oarg_96_din),
        .ap_fifo_oarg_96_write(ap_fifo_oarg_96_write),
        .m_axis_fifo_97_tlast(m_axis_fifo_97_tlast),
        .m_axis_fifo_97_tvalid(m_axis_fifo_97_tvalid),
        .m_axis_fifo_97_tkeep(m_axis_fifo_97_tkeep),
        .m_axis_fifo_97_tstrb(m_axis_fifo_97_tstrb),
        .m_axis_fifo_97_tdata(m_axis_fifo_97_tdata),
        .m_axis_fifo_97_tready(m_axis_fifo_97_tready),
        .ap_fifo_oarg_97_full_n(ap_fifo_oarg_97_full_n),
        .ap_fifo_oarg_97_din(ap_fifo_oarg_97_din),
        .ap_fifo_oarg_97_write(ap_fifo_oarg_97_write),
        .m_axis_fifo_98_tlast(m_axis_fifo_98_tlast),
        .m_axis_fifo_98_tvalid(m_axis_fifo_98_tvalid),
        .m_axis_fifo_98_tkeep(m_axis_fifo_98_tkeep),
        .m_axis_fifo_98_tstrb(m_axis_fifo_98_tstrb),
        .m_axis_fifo_98_tdata(m_axis_fifo_98_tdata),
        .m_axis_fifo_98_tready(m_axis_fifo_98_tready),
        .ap_fifo_oarg_98_full_n(ap_fifo_oarg_98_full_n),
        .ap_fifo_oarg_98_din(ap_fifo_oarg_98_din),
        .ap_fifo_oarg_98_write(ap_fifo_oarg_98_write),
        .m_axis_fifo_99_tlast(m_axis_fifo_99_tlast),
        .m_axis_fifo_99_tvalid(m_axis_fifo_99_tvalid),
        .m_axis_fifo_99_tkeep(m_axis_fifo_99_tkeep),
        .m_axis_fifo_99_tstrb(m_axis_fifo_99_tstrb),
        .m_axis_fifo_99_tdata(m_axis_fifo_99_tdata),
        .m_axis_fifo_99_tready(m_axis_fifo_99_tready),
        .ap_fifo_oarg_99_full_n(ap_fifo_oarg_99_full_n),
        .ap_fifo_oarg_99_din(ap_fifo_oarg_99_din),
        .ap_fifo_oarg_99_write(ap_fifo_oarg_99_write),
        .m_axis_fifo_100_tlast(m_axis_fifo_100_tlast),
        .m_axis_fifo_100_tvalid(m_axis_fifo_100_tvalid),
        .m_axis_fifo_100_tkeep(m_axis_fifo_100_tkeep),
        .m_axis_fifo_100_tstrb(m_axis_fifo_100_tstrb),
        .m_axis_fifo_100_tdata(m_axis_fifo_100_tdata),
        .m_axis_fifo_100_tready(m_axis_fifo_100_tready),
        .ap_fifo_oarg_100_full_n(ap_fifo_oarg_100_full_n),
        .ap_fifo_oarg_100_din(ap_fifo_oarg_100_din),
        .ap_fifo_oarg_100_write(ap_fifo_oarg_100_write),
        .m_axis_fifo_101_tlast(m_axis_fifo_101_tlast),
        .m_axis_fifo_101_tvalid(m_axis_fifo_101_tvalid),
        .m_axis_fifo_101_tkeep(m_axis_fifo_101_tkeep),
        .m_axis_fifo_101_tstrb(m_axis_fifo_101_tstrb),
        .m_axis_fifo_101_tdata(m_axis_fifo_101_tdata),
        .m_axis_fifo_101_tready(m_axis_fifo_101_tready),
        .ap_fifo_oarg_101_full_n(ap_fifo_oarg_101_full_n),
        .ap_fifo_oarg_101_din(ap_fifo_oarg_101_din),
        .ap_fifo_oarg_101_write(ap_fifo_oarg_101_write),
        .m_axis_fifo_102_tlast(m_axis_fifo_102_tlast),
        .m_axis_fifo_102_tvalid(m_axis_fifo_102_tvalid),
        .m_axis_fifo_102_tkeep(m_axis_fifo_102_tkeep),
        .m_axis_fifo_102_tstrb(m_axis_fifo_102_tstrb),
        .m_axis_fifo_102_tdata(m_axis_fifo_102_tdata),
        .m_axis_fifo_102_tready(m_axis_fifo_102_tready),
        .ap_fifo_oarg_102_full_n(ap_fifo_oarg_102_full_n),
        .ap_fifo_oarg_102_din(ap_fifo_oarg_102_din),
        .ap_fifo_oarg_102_write(ap_fifo_oarg_102_write),
        .m_axis_fifo_103_tlast(m_axis_fifo_103_tlast),
        .m_axis_fifo_103_tvalid(m_axis_fifo_103_tvalid),
        .m_axis_fifo_103_tkeep(m_axis_fifo_103_tkeep),
        .m_axis_fifo_103_tstrb(m_axis_fifo_103_tstrb),
        .m_axis_fifo_103_tdata(m_axis_fifo_103_tdata),
        .m_axis_fifo_103_tready(m_axis_fifo_103_tready),
        .ap_fifo_oarg_103_full_n(ap_fifo_oarg_103_full_n),
        .ap_fifo_oarg_103_din(ap_fifo_oarg_103_din),
        .ap_fifo_oarg_103_write(ap_fifo_oarg_103_write),
        .m_axis_fifo_104_tlast(m_axis_fifo_104_tlast),
        .m_axis_fifo_104_tvalid(m_axis_fifo_104_tvalid),
        .m_axis_fifo_104_tkeep(m_axis_fifo_104_tkeep),
        .m_axis_fifo_104_tstrb(m_axis_fifo_104_tstrb),
        .m_axis_fifo_104_tdata(m_axis_fifo_104_tdata),
        .m_axis_fifo_104_tready(m_axis_fifo_104_tready),
        .ap_fifo_oarg_104_full_n(ap_fifo_oarg_104_full_n),
        .ap_fifo_oarg_104_din(ap_fifo_oarg_104_din),
        .ap_fifo_oarg_104_write(ap_fifo_oarg_104_write),
        .m_axis_fifo_105_tlast(m_axis_fifo_105_tlast),
        .m_axis_fifo_105_tvalid(m_axis_fifo_105_tvalid),
        .m_axis_fifo_105_tkeep(m_axis_fifo_105_tkeep),
        .m_axis_fifo_105_tstrb(m_axis_fifo_105_tstrb),
        .m_axis_fifo_105_tdata(m_axis_fifo_105_tdata),
        .m_axis_fifo_105_tready(m_axis_fifo_105_tready),
        .ap_fifo_oarg_105_full_n(ap_fifo_oarg_105_full_n),
        .ap_fifo_oarg_105_din(ap_fifo_oarg_105_din),
        .ap_fifo_oarg_105_write(ap_fifo_oarg_105_write),
        .m_axis_fifo_106_tlast(m_axis_fifo_106_tlast),
        .m_axis_fifo_106_tvalid(m_axis_fifo_106_tvalid),
        .m_axis_fifo_106_tkeep(m_axis_fifo_106_tkeep),
        .m_axis_fifo_106_tstrb(m_axis_fifo_106_tstrb),
        .m_axis_fifo_106_tdata(m_axis_fifo_106_tdata),
        .m_axis_fifo_106_tready(m_axis_fifo_106_tready),
        .ap_fifo_oarg_106_full_n(ap_fifo_oarg_106_full_n),
        .ap_fifo_oarg_106_din(ap_fifo_oarg_106_din),
        .ap_fifo_oarg_106_write(ap_fifo_oarg_106_write),
        .m_axis_fifo_107_tlast(m_axis_fifo_107_tlast),
        .m_axis_fifo_107_tvalid(m_axis_fifo_107_tvalid),
        .m_axis_fifo_107_tkeep(m_axis_fifo_107_tkeep),
        .m_axis_fifo_107_tstrb(m_axis_fifo_107_tstrb),
        .m_axis_fifo_107_tdata(m_axis_fifo_107_tdata),
        .m_axis_fifo_107_tready(m_axis_fifo_107_tready),
        .ap_fifo_oarg_107_full_n(ap_fifo_oarg_107_full_n),
        .ap_fifo_oarg_107_din(ap_fifo_oarg_107_din),
        .ap_fifo_oarg_107_write(ap_fifo_oarg_107_write),
        .m_axis_fifo_108_tlast(m_axis_fifo_108_tlast),
        .m_axis_fifo_108_tvalid(m_axis_fifo_108_tvalid),
        .m_axis_fifo_108_tkeep(m_axis_fifo_108_tkeep),
        .m_axis_fifo_108_tstrb(m_axis_fifo_108_tstrb),
        .m_axis_fifo_108_tdata(m_axis_fifo_108_tdata),
        .m_axis_fifo_108_tready(m_axis_fifo_108_tready),
        .ap_fifo_oarg_108_full_n(ap_fifo_oarg_108_full_n),
        .ap_fifo_oarg_108_din(ap_fifo_oarg_108_din),
        .ap_fifo_oarg_108_write(ap_fifo_oarg_108_write),
        .m_axis_fifo_109_tlast(m_axis_fifo_109_tlast),
        .m_axis_fifo_109_tvalid(m_axis_fifo_109_tvalid),
        .m_axis_fifo_109_tkeep(m_axis_fifo_109_tkeep),
        .m_axis_fifo_109_tstrb(m_axis_fifo_109_tstrb),
        .m_axis_fifo_109_tdata(m_axis_fifo_109_tdata),
        .m_axis_fifo_109_tready(m_axis_fifo_109_tready),
        .ap_fifo_oarg_109_full_n(ap_fifo_oarg_109_full_n),
        .ap_fifo_oarg_109_din(ap_fifo_oarg_109_din),
        .ap_fifo_oarg_109_write(ap_fifo_oarg_109_write),
        .m_axis_fifo_110_tlast(m_axis_fifo_110_tlast),
        .m_axis_fifo_110_tvalid(m_axis_fifo_110_tvalid),
        .m_axis_fifo_110_tkeep(m_axis_fifo_110_tkeep),
        .m_axis_fifo_110_tstrb(m_axis_fifo_110_tstrb),
        .m_axis_fifo_110_tdata(m_axis_fifo_110_tdata),
        .m_axis_fifo_110_tready(m_axis_fifo_110_tready),
        .ap_fifo_oarg_110_full_n(ap_fifo_oarg_110_full_n),
        .ap_fifo_oarg_110_din(ap_fifo_oarg_110_din),
        .ap_fifo_oarg_110_write(ap_fifo_oarg_110_write),
        .m_axis_fifo_111_tlast(m_axis_fifo_111_tlast),
        .m_axis_fifo_111_tvalid(m_axis_fifo_111_tvalid),
        .m_axis_fifo_111_tkeep(m_axis_fifo_111_tkeep),
        .m_axis_fifo_111_tstrb(m_axis_fifo_111_tstrb),
        .m_axis_fifo_111_tdata(m_axis_fifo_111_tdata),
        .m_axis_fifo_111_tready(m_axis_fifo_111_tready),
        .ap_fifo_oarg_111_full_n(ap_fifo_oarg_111_full_n),
        .ap_fifo_oarg_111_din(ap_fifo_oarg_111_din),
        .ap_fifo_oarg_111_write(ap_fifo_oarg_111_write),
        .m_axis_fifo_112_tlast(m_axis_fifo_112_tlast),
        .m_axis_fifo_112_tvalid(m_axis_fifo_112_tvalid),
        .m_axis_fifo_112_tkeep(m_axis_fifo_112_tkeep),
        .m_axis_fifo_112_tstrb(m_axis_fifo_112_tstrb),
        .m_axis_fifo_112_tdata(m_axis_fifo_112_tdata),
        .m_axis_fifo_112_tready(m_axis_fifo_112_tready),
        .ap_fifo_oarg_112_full_n(ap_fifo_oarg_112_full_n),
        .ap_fifo_oarg_112_din(ap_fifo_oarg_112_din),
        .ap_fifo_oarg_112_write(ap_fifo_oarg_112_write),
        .m_axis_fifo_113_tlast(m_axis_fifo_113_tlast),
        .m_axis_fifo_113_tvalid(m_axis_fifo_113_tvalid),
        .m_axis_fifo_113_tkeep(m_axis_fifo_113_tkeep),
        .m_axis_fifo_113_tstrb(m_axis_fifo_113_tstrb),
        .m_axis_fifo_113_tdata(m_axis_fifo_113_tdata),
        .m_axis_fifo_113_tready(m_axis_fifo_113_tready),
        .ap_fifo_oarg_113_full_n(ap_fifo_oarg_113_full_n),
        .ap_fifo_oarg_113_din(ap_fifo_oarg_113_din),
        .ap_fifo_oarg_113_write(ap_fifo_oarg_113_write),
        .m_axis_fifo_114_tlast(m_axis_fifo_114_tlast),
        .m_axis_fifo_114_tvalid(m_axis_fifo_114_tvalid),
        .m_axis_fifo_114_tkeep(m_axis_fifo_114_tkeep),
        .m_axis_fifo_114_tstrb(m_axis_fifo_114_tstrb),
        .m_axis_fifo_114_tdata(m_axis_fifo_114_tdata),
        .m_axis_fifo_114_tready(m_axis_fifo_114_tready),
        .ap_fifo_oarg_114_full_n(ap_fifo_oarg_114_full_n),
        .ap_fifo_oarg_114_din(ap_fifo_oarg_114_din),
        .ap_fifo_oarg_114_write(ap_fifo_oarg_114_write),
        .m_axis_fifo_115_tlast(m_axis_fifo_115_tlast),
        .m_axis_fifo_115_tvalid(m_axis_fifo_115_tvalid),
        .m_axis_fifo_115_tkeep(m_axis_fifo_115_tkeep),
        .m_axis_fifo_115_tstrb(m_axis_fifo_115_tstrb),
        .m_axis_fifo_115_tdata(m_axis_fifo_115_tdata),
        .m_axis_fifo_115_tready(m_axis_fifo_115_tready),
        .ap_fifo_oarg_115_full_n(ap_fifo_oarg_115_full_n),
        .ap_fifo_oarg_115_din(ap_fifo_oarg_115_din),
        .ap_fifo_oarg_115_write(ap_fifo_oarg_115_write),
        .m_axis_fifo_116_tlast(m_axis_fifo_116_tlast),
        .m_axis_fifo_116_tvalid(m_axis_fifo_116_tvalid),
        .m_axis_fifo_116_tkeep(m_axis_fifo_116_tkeep),
        .m_axis_fifo_116_tstrb(m_axis_fifo_116_tstrb),
        .m_axis_fifo_116_tdata(m_axis_fifo_116_tdata),
        .m_axis_fifo_116_tready(m_axis_fifo_116_tready),
        .ap_fifo_oarg_116_full_n(ap_fifo_oarg_116_full_n),
        .ap_fifo_oarg_116_din(ap_fifo_oarg_116_din),
        .ap_fifo_oarg_116_write(ap_fifo_oarg_116_write),
        .m_axis_fifo_117_tlast(m_axis_fifo_117_tlast),
        .m_axis_fifo_117_tvalid(m_axis_fifo_117_tvalid),
        .m_axis_fifo_117_tkeep(m_axis_fifo_117_tkeep),
        .m_axis_fifo_117_tstrb(m_axis_fifo_117_tstrb),
        .m_axis_fifo_117_tdata(m_axis_fifo_117_tdata),
        .m_axis_fifo_117_tready(m_axis_fifo_117_tready),
        .ap_fifo_oarg_117_full_n(ap_fifo_oarg_117_full_n),
        .ap_fifo_oarg_117_din(ap_fifo_oarg_117_din),
        .ap_fifo_oarg_117_write(ap_fifo_oarg_117_write),
        .m_axis_fifo_118_tlast(m_axis_fifo_118_tlast),
        .m_axis_fifo_118_tvalid(m_axis_fifo_118_tvalid),
        .m_axis_fifo_118_tkeep(m_axis_fifo_118_tkeep),
        .m_axis_fifo_118_tstrb(m_axis_fifo_118_tstrb),
        .m_axis_fifo_118_tdata(m_axis_fifo_118_tdata),
        .m_axis_fifo_118_tready(m_axis_fifo_118_tready),
        .ap_fifo_oarg_118_full_n(ap_fifo_oarg_118_full_n),
        .ap_fifo_oarg_118_din(ap_fifo_oarg_118_din),
        .ap_fifo_oarg_118_write(ap_fifo_oarg_118_write),
        .m_axis_fifo_119_tlast(m_axis_fifo_119_tlast),
        .m_axis_fifo_119_tvalid(m_axis_fifo_119_tvalid),
        .m_axis_fifo_119_tkeep(m_axis_fifo_119_tkeep),
        .m_axis_fifo_119_tstrb(m_axis_fifo_119_tstrb),
        .m_axis_fifo_119_tdata(m_axis_fifo_119_tdata),
        .m_axis_fifo_119_tready(m_axis_fifo_119_tready),
        .ap_fifo_oarg_119_full_n(ap_fifo_oarg_119_full_n),
        .ap_fifo_oarg_119_din(ap_fifo_oarg_119_din),
        .ap_fifo_oarg_119_write(ap_fifo_oarg_119_write),
        .m_axis_fifo_120_tlast(m_axis_fifo_120_tlast),
        .m_axis_fifo_120_tvalid(m_axis_fifo_120_tvalid),
        .m_axis_fifo_120_tkeep(m_axis_fifo_120_tkeep),
        .m_axis_fifo_120_tstrb(m_axis_fifo_120_tstrb),
        .m_axis_fifo_120_tdata(m_axis_fifo_120_tdata),
        .m_axis_fifo_120_tready(m_axis_fifo_120_tready),
        .ap_fifo_oarg_120_full_n(ap_fifo_oarg_120_full_n),
        .ap_fifo_oarg_120_din(ap_fifo_oarg_120_din),
        .ap_fifo_oarg_120_write(ap_fifo_oarg_120_write),
        .m_axis_fifo_121_tlast(m_axis_fifo_121_tlast),
        .m_axis_fifo_121_tvalid(m_axis_fifo_121_tvalid),
        .m_axis_fifo_121_tkeep(m_axis_fifo_121_tkeep),
        .m_axis_fifo_121_tstrb(m_axis_fifo_121_tstrb),
        .m_axis_fifo_121_tdata(m_axis_fifo_121_tdata),
        .m_axis_fifo_121_tready(m_axis_fifo_121_tready),
        .ap_fifo_oarg_121_full_n(ap_fifo_oarg_121_full_n),
        .ap_fifo_oarg_121_din(ap_fifo_oarg_121_din),
        .ap_fifo_oarg_121_write(ap_fifo_oarg_121_write),
        .m_axis_fifo_122_tlast(m_axis_fifo_122_tlast),
        .m_axis_fifo_122_tvalid(m_axis_fifo_122_tvalid),
        .m_axis_fifo_122_tkeep(m_axis_fifo_122_tkeep),
        .m_axis_fifo_122_tstrb(m_axis_fifo_122_tstrb),
        .m_axis_fifo_122_tdata(m_axis_fifo_122_tdata),
        .m_axis_fifo_122_tready(m_axis_fifo_122_tready),
        .ap_fifo_oarg_122_full_n(ap_fifo_oarg_122_full_n),
        .ap_fifo_oarg_122_din(ap_fifo_oarg_122_din),
        .ap_fifo_oarg_122_write(ap_fifo_oarg_122_write),
        .m_axis_fifo_123_tlast(m_axis_fifo_123_tlast),
        .m_axis_fifo_123_tvalid(m_axis_fifo_123_tvalid),
        .m_axis_fifo_123_tkeep(m_axis_fifo_123_tkeep),
        .m_axis_fifo_123_tstrb(m_axis_fifo_123_tstrb),
        .m_axis_fifo_123_tdata(m_axis_fifo_123_tdata),
        .m_axis_fifo_123_tready(m_axis_fifo_123_tready),
        .ap_fifo_oarg_123_full_n(ap_fifo_oarg_123_full_n),
        .ap_fifo_oarg_123_din(ap_fifo_oarg_123_din),
        .ap_fifo_oarg_123_write(ap_fifo_oarg_123_write),
        .m_axis_fifo_124_tlast(m_axis_fifo_124_tlast),
        .m_axis_fifo_124_tvalid(m_axis_fifo_124_tvalid),
        .m_axis_fifo_124_tkeep(m_axis_fifo_124_tkeep),
        .m_axis_fifo_124_tstrb(m_axis_fifo_124_tstrb),
        .m_axis_fifo_124_tdata(m_axis_fifo_124_tdata),
        .m_axis_fifo_124_tready(m_axis_fifo_124_tready),
        .ap_fifo_oarg_124_full_n(ap_fifo_oarg_124_full_n),
        .ap_fifo_oarg_124_din(ap_fifo_oarg_124_din),
        .ap_fifo_oarg_124_write(ap_fifo_oarg_124_write),
        .m_axis_fifo_125_tlast(m_axis_fifo_125_tlast),
        .m_axis_fifo_125_tvalid(m_axis_fifo_125_tvalid),
        .m_axis_fifo_125_tkeep(m_axis_fifo_125_tkeep),
        .m_axis_fifo_125_tstrb(m_axis_fifo_125_tstrb),
        .m_axis_fifo_125_tdata(m_axis_fifo_125_tdata),
        .m_axis_fifo_125_tready(m_axis_fifo_125_tready),
        .ap_fifo_oarg_125_full_n(ap_fifo_oarg_125_full_n),
        .ap_fifo_oarg_125_din(ap_fifo_oarg_125_din),
        .ap_fifo_oarg_125_write(ap_fifo_oarg_125_write),
        .m_axis_fifo_126_tlast(m_axis_fifo_126_tlast),
        .m_axis_fifo_126_tvalid(m_axis_fifo_126_tvalid),
        .m_axis_fifo_126_tkeep(m_axis_fifo_126_tkeep),
        .m_axis_fifo_126_tstrb(m_axis_fifo_126_tstrb),
        .m_axis_fifo_126_tdata(m_axis_fifo_126_tdata),
        .m_axis_fifo_126_tready(m_axis_fifo_126_tready),
        .ap_fifo_oarg_126_full_n(ap_fifo_oarg_126_full_n),
        .ap_fifo_oarg_126_din(ap_fifo_oarg_126_din),
        .ap_fifo_oarg_126_write(ap_fifo_oarg_126_write),
        .m_axis_fifo_127_tlast(m_axis_fifo_127_tlast),
        .m_axis_fifo_127_tvalid(m_axis_fifo_127_tvalid),
        .m_axis_fifo_127_tkeep(m_axis_fifo_127_tkeep),
        .m_axis_fifo_127_tstrb(m_axis_fifo_127_tstrb),
        .m_axis_fifo_127_tdata(m_axis_fifo_127_tdata),
        .m_axis_fifo_127_tready(m_axis_fifo_127_tready),
        .ap_fifo_oarg_127_full_n(ap_fifo_oarg_127_full_n),
        .ap_fifo_oarg_127_din(ap_fifo_oarg_127_din),
        .ap_fifo_oarg_127_write(ap_fifo_oarg_127_write)
    );
    
    in_bram_args #(
        .C_NUM_INPUT_BRAMs(C_NUM_INPUT_BRAMs),
        .C_INPUT_BRAM_0_PORTS(C_INPUT_BRAM_0_PORTS),
        .C_INPUT_BRAM_1_PORTS(C_INPUT_BRAM_1_PORTS),
        .C_INPUT_BRAM_2_PORTS(C_INPUT_BRAM_2_PORTS),
        .C_INPUT_BRAM_3_PORTS(C_INPUT_BRAM_3_PORTS),
        .C_INPUT_BRAM_4_PORTS(C_INPUT_BRAM_4_PORTS),
        .C_INPUT_BRAM_5_PORTS(C_INPUT_BRAM_5_PORTS),
        .C_INPUT_BRAM_6_PORTS(C_INPUT_BRAM_6_PORTS),
        .C_INPUT_BRAM_7_PORTS(C_INPUT_BRAM_7_PORTS),
        .C_INPUT_BRAM_8_PORTS(C_INPUT_BRAM_8_PORTS),
        .C_INPUT_BRAM_9_PORTS(C_INPUT_BRAM_9_PORTS),
        .C_INPUT_BRAM_10_PORTS(C_INPUT_BRAM_10_PORTS),
        .C_INPUT_BRAM_11_PORTS(C_INPUT_BRAM_11_PORTS),
        .C_INPUT_BRAM_12_PORTS(C_INPUT_BRAM_12_PORTS),
        .C_INPUT_BRAM_13_PORTS(C_INPUT_BRAM_13_PORTS),
        .C_INPUT_BRAM_14_PORTS(C_INPUT_BRAM_14_PORTS),
        .C_INPUT_BRAM_15_PORTS(C_INPUT_BRAM_15_PORTS),
        .C_INPUT_BRAM_16_PORTS(C_INPUT_BRAM_16_PORTS),
        .C_INPUT_BRAM_17_PORTS(C_INPUT_BRAM_17_PORTS),
        .C_INPUT_BRAM_18_PORTS(C_INPUT_BRAM_18_PORTS),
        .C_INPUT_BRAM_19_PORTS(C_INPUT_BRAM_19_PORTS),
        .C_INPUT_BRAM_20_PORTS(C_INPUT_BRAM_20_PORTS),
        .C_INPUT_BRAM_21_PORTS(C_INPUT_BRAM_21_PORTS),
        .C_INPUT_BRAM_22_PORTS(C_INPUT_BRAM_22_PORTS),
        .C_INPUT_BRAM_23_PORTS(C_INPUT_BRAM_23_PORTS),
        .C_INPUT_BRAM_24_PORTS(C_INPUT_BRAM_24_PORTS),
        .C_INPUT_BRAM_25_PORTS(C_INPUT_BRAM_25_PORTS),
        .C_INPUT_BRAM_26_PORTS(C_INPUT_BRAM_26_PORTS),
        .C_INPUT_BRAM_27_PORTS(C_INPUT_BRAM_27_PORTS),
        .C_INPUT_BRAM_28_PORTS(C_INPUT_BRAM_28_PORTS),
        .C_INPUT_BRAM_29_PORTS(C_INPUT_BRAM_29_PORTS),
        .C_INPUT_BRAM_30_PORTS(C_INPUT_BRAM_30_PORTS),
        .C_INPUT_BRAM_31_PORTS(C_INPUT_BRAM_31_PORTS),
        .C_INPUT_BRAM_32_PORTS(C_INPUT_BRAM_32_PORTS),
        .C_INPUT_BRAM_33_PORTS(C_INPUT_BRAM_33_PORTS),
        .C_INPUT_BRAM_34_PORTS(C_INPUT_BRAM_34_PORTS),
        .C_INPUT_BRAM_35_PORTS(C_INPUT_BRAM_35_PORTS),
        .C_INPUT_BRAM_36_PORTS(C_INPUT_BRAM_36_PORTS),
        .C_INPUT_BRAM_37_PORTS(C_INPUT_BRAM_37_PORTS),
        .C_INPUT_BRAM_38_PORTS(C_INPUT_BRAM_38_PORTS),
        .C_INPUT_BRAM_39_PORTS(C_INPUT_BRAM_39_PORTS),
        .C_INPUT_BRAM_40_PORTS(C_INPUT_BRAM_40_PORTS),
        .C_INPUT_BRAM_41_PORTS(C_INPUT_BRAM_41_PORTS),
        .C_INPUT_BRAM_42_PORTS(C_INPUT_BRAM_42_PORTS),
        .C_INPUT_BRAM_43_PORTS(C_INPUT_BRAM_43_PORTS),
        .C_INPUT_BRAM_44_PORTS(C_INPUT_BRAM_44_PORTS),
        .C_INPUT_BRAM_45_PORTS(C_INPUT_BRAM_45_PORTS),
        .C_INPUT_BRAM_46_PORTS(C_INPUT_BRAM_46_PORTS),
        .C_INPUT_BRAM_47_PORTS(C_INPUT_BRAM_47_PORTS),
        .C_INPUT_BRAM_48_PORTS(C_INPUT_BRAM_48_PORTS),
        .C_INPUT_BRAM_49_PORTS(C_INPUT_BRAM_49_PORTS),
        .C_INPUT_BRAM_50_PORTS(C_INPUT_BRAM_50_PORTS),
        .C_INPUT_BRAM_51_PORTS(C_INPUT_BRAM_51_PORTS),
        .C_INPUT_BRAM_52_PORTS(C_INPUT_BRAM_52_PORTS),
        .C_INPUT_BRAM_53_PORTS(C_INPUT_BRAM_53_PORTS),
        .C_INPUT_BRAM_54_PORTS(C_INPUT_BRAM_54_PORTS),
        .C_INPUT_BRAM_55_PORTS(C_INPUT_BRAM_55_PORTS),
        .C_INPUT_BRAM_56_PORTS(C_INPUT_BRAM_56_PORTS),
        .C_INPUT_BRAM_57_PORTS(C_INPUT_BRAM_57_PORTS),
        .C_INPUT_BRAM_58_PORTS(C_INPUT_BRAM_58_PORTS),
        .C_INPUT_BRAM_59_PORTS(C_INPUT_BRAM_59_PORTS),
        .C_INPUT_BRAM_60_PORTS(C_INPUT_BRAM_60_PORTS),
        .C_INPUT_BRAM_61_PORTS(C_INPUT_BRAM_61_PORTS),
        .C_INPUT_BRAM_62_PORTS(C_INPUT_BRAM_62_PORTS),
        .C_INPUT_BRAM_63_PORTS(C_INPUT_BRAM_63_PORTS),
        .C_INPUT_BRAM_64_PORTS(C_INPUT_BRAM_64_PORTS),
        .C_INPUT_BRAM_65_PORTS(C_INPUT_BRAM_65_PORTS),
        .C_INPUT_BRAM_66_PORTS(C_INPUT_BRAM_66_PORTS),
        .C_INPUT_BRAM_67_PORTS(C_INPUT_BRAM_67_PORTS),
        .C_INPUT_BRAM_68_PORTS(C_INPUT_BRAM_68_PORTS),
        .C_INPUT_BRAM_69_PORTS(C_INPUT_BRAM_69_PORTS),
        .C_INPUT_BRAM_70_PORTS(C_INPUT_BRAM_70_PORTS),
        .C_INPUT_BRAM_71_PORTS(C_INPUT_BRAM_71_PORTS),
        .C_INPUT_BRAM_72_PORTS(C_INPUT_BRAM_72_PORTS),
        .C_INPUT_BRAM_73_PORTS(C_INPUT_BRAM_73_PORTS),
        .C_INPUT_BRAM_74_PORTS(C_INPUT_BRAM_74_PORTS),
        .C_INPUT_BRAM_75_PORTS(C_INPUT_BRAM_75_PORTS),
        .C_INPUT_BRAM_76_PORTS(C_INPUT_BRAM_76_PORTS),
        .C_INPUT_BRAM_77_PORTS(C_INPUT_BRAM_77_PORTS),
        .C_INPUT_BRAM_78_PORTS(C_INPUT_BRAM_78_PORTS),
        .C_INPUT_BRAM_79_PORTS(C_INPUT_BRAM_79_PORTS),
        .C_INPUT_BRAM_80_PORTS(C_INPUT_BRAM_80_PORTS),
        .C_INPUT_BRAM_81_PORTS(C_INPUT_BRAM_81_PORTS),
        .C_INPUT_BRAM_82_PORTS(C_INPUT_BRAM_82_PORTS),
        .C_INPUT_BRAM_83_PORTS(C_INPUT_BRAM_83_PORTS),
        .C_INPUT_BRAM_84_PORTS(C_INPUT_BRAM_84_PORTS),
        .C_INPUT_BRAM_85_PORTS(C_INPUT_BRAM_85_PORTS),
        .C_INPUT_BRAM_86_PORTS(C_INPUT_BRAM_86_PORTS),
        .C_INPUT_BRAM_87_PORTS(C_INPUT_BRAM_87_PORTS),
        .C_INPUT_BRAM_88_PORTS(C_INPUT_BRAM_88_PORTS),
        .C_INPUT_BRAM_89_PORTS(C_INPUT_BRAM_89_PORTS),
        .C_INPUT_BRAM_90_PORTS(C_INPUT_BRAM_90_PORTS),
        .C_INPUT_BRAM_91_PORTS(C_INPUT_BRAM_91_PORTS),
        .C_INPUT_BRAM_92_PORTS(C_INPUT_BRAM_92_PORTS),
        .C_INPUT_BRAM_93_PORTS(C_INPUT_BRAM_93_PORTS),
        .C_INPUT_BRAM_94_PORTS(C_INPUT_BRAM_94_PORTS),
        .C_INPUT_BRAM_95_PORTS(C_INPUT_BRAM_95_PORTS),
        .C_INPUT_BRAM_96_PORTS(C_INPUT_BRAM_96_PORTS),
        .C_INPUT_BRAM_97_PORTS(C_INPUT_BRAM_97_PORTS),
        .C_INPUT_BRAM_98_PORTS(C_INPUT_BRAM_98_PORTS),
        .C_INPUT_BRAM_99_PORTS(C_INPUT_BRAM_99_PORTS),
        .C_INPUT_BRAM_100_PORTS(C_INPUT_BRAM_100_PORTS),
        .C_INPUT_BRAM_101_PORTS(C_INPUT_BRAM_101_PORTS),
        .C_INPUT_BRAM_102_PORTS(C_INPUT_BRAM_102_PORTS),
        .C_INPUT_BRAM_103_PORTS(C_INPUT_BRAM_103_PORTS),
        .C_INPUT_BRAM_104_PORTS(C_INPUT_BRAM_104_PORTS),
        .C_INPUT_BRAM_105_PORTS(C_INPUT_BRAM_105_PORTS),
        .C_INPUT_BRAM_106_PORTS(C_INPUT_BRAM_106_PORTS),
        .C_INPUT_BRAM_107_PORTS(C_INPUT_BRAM_107_PORTS),
        .C_INPUT_BRAM_108_PORTS(C_INPUT_BRAM_108_PORTS),
        .C_INPUT_BRAM_109_PORTS(C_INPUT_BRAM_109_PORTS),
        .C_INPUT_BRAM_110_PORTS(C_INPUT_BRAM_110_PORTS),
        .C_INPUT_BRAM_111_PORTS(C_INPUT_BRAM_111_PORTS),
        .C_INPUT_BRAM_112_PORTS(C_INPUT_BRAM_112_PORTS),
        .C_INPUT_BRAM_113_PORTS(C_INPUT_BRAM_113_PORTS),
        .C_INPUT_BRAM_114_PORTS(C_INPUT_BRAM_114_PORTS),
        .C_INPUT_BRAM_115_PORTS(C_INPUT_BRAM_115_PORTS),
        .C_INPUT_BRAM_116_PORTS(C_INPUT_BRAM_116_PORTS),
        .C_INPUT_BRAM_117_PORTS(C_INPUT_BRAM_117_PORTS),
        .C_INPUT_BRAM_118_PORTS(C_INPUT_BRAM_118_PORTS),
        .C_INPUT_BRAM_119_PORTS(C_INPUT_BRAM_119_PORTS),
        .C_INPUT_BRAM_120_PORTS(C_INPUT_BRAM_120_PORTS),
        .C_INPUT_BRAM_121_PORTS(C_INPUT_BRAM_121_PORTS),
        .C_INPUT_BRAM_122_PORTS(C_INPUT_BRAM_122_PORTS),
        .C_INPUT_BRAM_123_PORTS(C_INPUT_BRAM_123_PORTS),
        .C_INPUT_BRAM_124_PORTS(C_INPUT_BRAM_124_PORTS),
        .C_INPUT_BRAM_125_PORTS(C_INPUT_BRAM_125_PORTS),
        .C_INPUT_BRAM_126_PORTS(C_INPUT_BRAM_126_PORTS),
        .C_INPUT_BRAM_127_PORTS(C_INPUT_BRAM_127_PORTS),
        .C_INPUT_BRAM_0_WIDTH(C_INPUT_BRAM_0_WIDTH),
        .C_INPUT_BRAM_1_WIDTH(C_INPUT_BRAM_1_WIDTH),
        .C_INPUT_BRAM_2_WIDTH(C_INPUT_BRAM_2_WIDTH),
        .C_INPUT_BRAM_3_WIDTH(C_INPUT_BRAM_3_WIDTH),
        .C_INPUT_BRAM_4_WIDTH(C_INPUT_BRAM_4_WIDTH),
        .C_INPUT_BRAM_5_WIDTH(C_INPUT_BRAM_5_WIDTH),
        .C_INPUT_BRAM_6_WIDTH(C_INPUT_BRAM_6_WIDTH),
        .C_INPUT_BRAM_7_WIDTH(C_INPUT_BRAM_7_WIDTH),
        .C_INPUT_BRAM_8_WIDTH(C_INPUT_BRAM_8_WIDTH),
        .C_INPUT_BRAM_9_WIDTH(C_INPUT_BRAM_9_WIDTH),
        .C_INPUT_BRAM_10_WIDTH(C_INPUT_BRAM_10_WIDTH),
        .C_INPUT_BRAM_11_WIDTH(C_INPUT_BRAM_11_WIDTH),
        .C_INPUT_BRAM_12_WIDTH(C_INPUT_BRAM_12_WIDTH),
        .C_INPUT_BRAM_13_WIDTH(C_INPUT_BRAM_13_WIDTH),
        .C_INPUT_BRAM_14_WIDTH(C_INPUT_BRAM_14_WIDTH),
        .C_INPUT_BRAM_15_WIDTH(C_INPUT_BRAM_15_WIDTH),
        .C_INPUT_BRAM_16_WIDTH(C_INPUT_BRAM_16_WIDTH),
        .C_INPUT_BRAM_17_WIDTH(C_INPUT_BRAM_17_WIDTH),
        .C_INPUT_BRAM_18_WIDTH(C_INPUT_BRAM_18_WIDTH),
        .C_INPUT_BRAM_19_WIDTH(C_INPUT_BRAM_19_WIDTH),
        .C_INPUT_BRAM_20_WIDTH(C_INPUT_BRAM_20_WIDTH),
        .C_INPUT_BRAM_21_WIDTH(C_INPUT_BRAM_21_WIDTH),
        .C_INPUT_BRAM_22_WIDTH(C_INPUT_BRAM_22_WIDTH),
        .C_INPUT_BRAM_23_WIDTH(C_INPUT_BRAM_23_WIDTH),
        .C_INPUT_BRAM_24_WIDTH(C_INPUT_BRAM_24_WIDTH),
        .C_INPUT_BRAM_25_WIDTH(C_INPUT_BRAM_25_WIDTH),
        .C_INPUT_BRAM_26_WIDTH(C_INPUT_BRAM_26_WIDTH),
        .C_INPUT_BRAM_27_WIDTH(C_INPUT_BRAM_27_WIDTH),
        .C_INPUT_BRAM_28_WIDTH(C_INPUT_BRAM_28_WIDTH),
        .C_INPUT_BRAM_29_WIDTH(C_INPUT_BRAM_29_WIDTH),
        .C_INPUT_BRAM_30_WIDTH(C_INPUT_BRAM_30_WIDTH),
        .C_INPUT_BRAM_31_WIDTH(C_INPUT_BRAM_31_WIDTH),
        .C_INPUT_BRAM_32_WIDTH(C_INPUT_BRAM_32_WIDTH),
        .C_INPUT_BRAM_33_WIDTH(C_INPUT_BRAM_33_WIDTH),
        .C_INPUT_BRAM_34_WIDTH(C_INPUT_BRAM_34_WIDTH),
        .C_INPUT_BRAM_35_WIDTH(C_INPUT_BRAM_35_WIDTH),
        .C_INPUT_BRAM_36_WIDTH(C_INPUT_BRAM_36_WIDTH),
        .C_INPUT_BRAM_37_WIDTH(C_INPUT_BRAM_37_WIDTH),
        .C_INPUT_BRAM_38_WIDTH(C_INPUT_BRAM_38_WIDTH),
        .C_INPUT_BRAM_39_WIDTH(C_INPUT_BRAM_39_WIDTH),
        .C_INPUT_BRAM_40_WIDTH(C_INPUT_BRAM_40_WIDTH),
        .C_INPUT_BRAM_41_WIDTH(C_INPUT_BRAM_41_WIDTH),
        .C_INPUT_BRAM_42_WIDTH(C_INPUT_BRAM_42_WIDTH),
        .C_INPUT_BRAM_43_WIDTH(C_INPUT_BRAM_43_WIDTH),
        .C_INPUT_BRAM_44_WIDTH(C_INPUT_BRAM_44_WIDTH),
        .C_INPUT_BRAM_45_WIDTH(C_INPUT_BRAM_45_WIDTH),
        .C_INPUT_BRAM_46_WIDTH(C_INPUT_BRAM_46_WIDTH),
        .C_INPUT_BRAM_47_WIDTH(C_INPUT_BRAM_47_WIDTH),
        .C_INPUT_BRAM_48_WIDTH(C_INPUT_BRAM_48_WIDTH),
        .C_INPUT_BRAM_49_WIDTH(C_INPUT_BRAM_49_WIDTH),
        .C_INPUT_BRAM_50_WIDTH(C_INPUT_BRAM_50_WIDTH),
        .C_INPUT_BRAM_51_WIDTH(C_INPUT_BRAM_51_WIDTH),
        .C_INPUT_BRAM_52_WIDTH(C_INPUT_BRAM_52_WIDTH),
        .C_INPUT_BRAM_53_WIDTH(C_INPUT_BRAM_53_WIDTH),
        .C_INPUT_BRAM_54_WIDTH(C_INPUT_BRAM_54_WIDTH),
        .C_INPUT_BRAM_55_WIDTH(C_INPUT_BRAM_55_WIDTH),
        .C_INPUT_BRAM_56_WIDTH(C_INPUT_BRAM_56_WIDTH),
        .C_INPUT_BRAM_57_WIDTH(C_INPUT_BRAM_57_WIDTH),
        .C_INPUT_BRAM_58_WIDTH(C_INPUT_BRAM_58_WIDTH),
        .C_INPUT_BRAM_59_WIDTH(C_INPUT_BRAM_59_WIDTH),
        .C_INPUT_BRAM_60_WIDTH(C_INPUT_BRAM_60_WIDTH),
        .C_INPUT_BRAM_61_WIDTH(C_INPUT_BRAM_61_WIDTH),
        .C_INPUT_BRAM_62_WIDTH(C_INPUT_BRAM_62_WIDTH),
        .C_INPUT_BRAM_63_WIDTH(C_INPUT_BRAM_63_WIDTH),
        .C_INPUT_BRAM_64_WIDTH(C_INPUT_BRAM_64_WIDTH),
        .C_INPUT_BRAM_65_WIDTH(C_INPUT_BRAM_65_WIDTH),
        .C_INPUT_BRAM_66_WIDTH(C_INPUT_BRAM_66_WIDTH),
        .C_INPUT_BRAM_67_WIDTH(C_INPUT_BRAM_67_WIDTH),
        .C_INPUT_BRAM_68_WIDTH(C_INPUT_BRAM_68_WIDTH),
        .C_INPUT_BRAM_69_WIDTH(C_INPUT_BRAM_69_WIDTH),
        .C_INPUT_BRAM_70_WIDTH(C_INPUT_BRAM_70_WIDTH),
        .C_INPUT_BRAM_71_WIDTH(C_INPUT_BRAM_71_WIDTH),
        .C_INPUT_BRAM_72_WIDTH(C_INPUT_BRAM_72_WIDTH),
        .C_INPUT_BRAM_73_WIDTH(C_INPUT_BRAM_73_WIDTH),
        .C_INPUT_BRAM_74_WIDTH(C_INPUT_BRAM_74_WIDTH),
        .C_INPUT_BRAM_75_WIDTH(C_INPUT_BRAM_75_WIDTH),
        .C_INPUT_BRAM_76_WIDTH(C_INPUT_BRAM_76_WIDTH),
        .C_INPUT_BRAM_77_WIDTH(C_INPUT_BRAM_77_WIDTH),
        .C_INPUT_BRAM_78_WIDTH(C_INPUT_BRAM_78_WIDTH),
        .C_INPUT_BRAM_79_WIDTH(C_INPUT_BRAM_79_WIDTH),
        .C_INPUT_BRAM_80_WIDTH(C_INPUT_BRAM_80_WIDTH),
        .C_INPUT_BRAM_81_WIDTH(C_INPUT_BRAM_81_WIDTH),
        .C_INPUT_BRAM_82_WIDTH(C_INPUT_BRAM_82_WIDTH),
        .C_INPUT_BRAM_83_WIDTH(C_INPUT_BRAM_83_WIDTH),
        .C_INPUT_BRAM_84_WIDTH(C_INPUT_BRAM_84_WIDTH),
        .C_INPUT_BRAM_85_WIDTH(C_INPUT_BRAM_85_WIDTH),
        .C_INPUT_BRAM_86_WIDTH(C_INPUT_BRAM_86_WIDTH),
        .C_INPUT_BRAM_87_WIDTH(C_INPUT_BRAM_87_WIDTH),
        .C_INPUT_BRAM_88_WIDTH(C_INPUT_BRAM_88_WIDTH),
        .C_INPUT_BRAM_89_WIDTH(C_INPUT_BRAM_89_WIDTH),
        .C_INPUT_BRAM_90_WIDTH(C_INPUT_BRAM_90_WIDTH),
        .C_INPUT_BRAM_91_WIDTH(C_INPUT_BRAM_91_WIDTH),
        .C_INPUT_BRAM_92_WIDTH(C_INPUT_BRAM_92_WIDTH),
        .C_INPUT_BRAM_93_WIDTH(C_INPUT_BRAM_93_WIDTH),
        .C_INPUT_BRAM_94_WIDTH(C_INPUT_BRAM_94_WIDTH),
        .C_INPUT_BRAM_95_WIDTH(C_INPUT_BRAM_95_WIDTH),
        .C_INPUT_BRAM_96_WIDTH(C_INPUT_BRAM_96_WIDTH),
        .C_INPUT_BRAM_97_WIDTH(C_INPUT_BRAM_97_WIDTH),
        .C_INPUT_BRAM_98_WIDTH(C_INPUT_BRAM_98_WIDTH),
        .C_INPUT_BRAM_99_WIDTH(C_INPUT_BRAM_99_WIDTH),
        .C_INPUT_BRAM_100_WIDTH(C_INPUT_BRAM_100_WIDTH),
        .C_INPUT_BRAM_101_WIDTH(C_INPUT_BRAM_101_WIDTH),
        .C_INPUT_BRAM_102_WIDTH(C_INPUT_BRAM_102_WIDTH),
        .C_INPUT_BRAM_103_WIDTH(C_INPUT_BRAM_103_WIDTH),
        .C_INPUT_BRAM_104_WIDTH(C_INPUT_BRAM_104_WIDTH),
        .C_INPUT_BRAM_105_WIDTH(C_INPUT_BRAM_105_WIDTH),
        .C_INPUT_BRAM_106_WIDTH(C_INPUT_BRAM_106_WIDTH),
        .C_INPUT_BRAM_107_WIDTH(C_INPUT_BRAM_107_WIDTH),
        .C_INPUT_BRAM_108_WIDTH(C_INPUT_BRAM_108_WIDTH),
        .C_INPUT_BRAM_109_WIDTH(C_INPUT_BRAM_109_WIDTH),
        .C_INPUT_BRAM_110_WIDTH(C_INPUT_BRAM_110_WIDTH),
        .C_INPUT_BRAM_111_WIDTH(C_INPUT_BRAM_111_WIDTH),
        .C_INPUT_BRAM_112_WIDTH(C_INPUT_BRAM_112_WIDTH),
        .C_INPUT_BRAM_113_WIDTH(C_INPUT_BRAM_113_WIDTH),
        .C_INPUT_BRAM_114_WIDTH(C_INPUT_BRAM_114_WIDTH),
        .C_INPUT_BRAM_115_WIDTH(C_INPUT_BRAM_115_WIDTH),
        .C_INPUT_BRAM_116_WIDTH(C_INPUT_BRAM_116_WIDTH),
        .C_INPUT_BRAM_117_WIDTH(C_INPUT_BRAM_117_WIDTH),
        .C_INPUT_BRAM_118_WIDTH(C_INPUT_BRAM_118_WIDTH),
        .C_INPUT_BRAM_119_WIDTH(C_INPUT_BRAM_119_WIDTH),
        .C_INPUT_BRAM_120_WIDTH(C_INPUT_BRAM_120_WIDTH),
        .C_INPUT_BRAM_121_WIDTH(C_INPUT_BRAM_121_WIDTH),
        .C_INPUT_BRAM_122_WIDTH(C_INPUT_BRAM_122_WIDTH),
        .C_INPUT_BRAM_123_WIDTH(C_INPUT_BRAM_123_WIDTH),
        .C_INPUT_BRAM_124_WIDTH(C_INPUT_BRAM_124_WIDTH),
        .C_INPUT_BRAM_125_WIDTH(C_INPUT_BRAM_125_WIDTH),
        .C_INPUT_BRAM_126_WIDTH(C_INPUT_BRAM_126_WIDTH),
        .C_INPUT_BRAM_127_WIDTH(C_INPUT_BRAM_127_WIDTH),
        .C_INPUT_BRAM_0_DEPTH(C_INPUT_BRAM_0_DEPTH),
        .C_INPUT_BRAM_1_DEPTH(C_INPUT_BRAM_1_DEPTH),
        .C_INPUT_BRAM_2_DEPTH(C_INPUT_BRAM_2_DEPTH),
        .C_INPUT_BRAM_3_DEPTH(C_INPUT_BRAM_3_DEPTH),
        .C_INPUT_BRAM_4_DEPTH(C_INPUT_BRAM_4_DEPTH),
        .C_INPUT_BRAM_5_DEPTH(C_INPUT_BRAM_5_DEPTH),
        .C_INPUT_BRAM_6_DEPTH(C_INPUT_BRAM_6_DEPTH),
        .C_INPUT_BRAM_7_DEPTH(C_INPUT_BRAM_7_DEPTH),
        .C_INPUT_BRAM_8_DEPTH(C_INPUT_BRAM_8_DEPTH),
        .C_INPUT_BRAM_9_DEPTH(C_INPUT_BRAM_9_DEPTH),
        .C_INPUT_BRAM_10_DEPTH(C_INPUT_BRAM_10_DEPTH),
        .C_INPUT_BRAM_11_DEPTH(C_INPUT_BRAM_11_DEPTH),
        .C_INPUT_BRAM_12_DEPTH(C_INPUT_BRAM_12_DEPTH),
        .C_INPUT_BRAM_13_DEPTH(C_INPUT_BRAM_13_DEPTH),
        .C_INPUT_BRAM_14_DEPTH(C_INPUT_BRAM_14_DEPTH),
        .C_INPUT_BRAM_15_DEPTH(C_INPUT_BRAM_15_DEPTH),
        .C_INPUT_BRAM_16_DEPTH(C_INPUT_BRAM_16_DEPTH),
        .C_INPUT_BRAM_17_DEPTH(C_INPUT_BRAM_17_DEPTH),
        .C_INPUT_BRAM_18_DEPTH(C_INPUT_BRAM_18_DEPTH),
        .C_INPUT_BRAM_19_DEPTH(C_INPUT_BRAM_19_DEPTH),
        .C_INPUT_BRAM_20_DEPTH(C_INPUT_BRAM_20_DEPTH),
        .C_INPUT_BRAM_21_DEPTH(C_INPUT_BRAM_21_DEPTH),
        .C_INPUT_BRAM_22_DEPTH(C_INPUT_BRAM_22_DEPTH),
        .C_INPUT_BRAM_23_DEPTH(C_INPUT_BRAM_23_DEPTH),
        .C_INPUT_BRAM_24_DEPTH(C_INPUT_BRAM_24_DEPTH),
        .C_INPUT_BRAM_25_DEPTH(C_INPUT_BRAM_25_DEPTH),
        .C_INPUT_BRAM_26_DEPTH(C_INPUT_BRAM_26_DEPTH),
        .C_INPUT_BRAM_27_DEPTH(C_INPUT_BRAM_27_DEPTH),
        .C_INPUT_BRAM_28_DEPTH(C_INPUT_BRAM_28_DEPTH),
        .C_INPUT_BRAM_29_DEPTH(C_INPUT_BRAM_29_DEPTH),
        .C_INPUT_BRAM_30_DEPTH(C_INPUT_BRAM_30_DEPTH),
        .C_INPUT_BRAM_31_DEPTH(C_INPUT_BRAM_31_DEPTH),
        .C_INPUT_BRAM_32_DEPTH(C_INPUT_BRAM_32_DEPTH),
        .C_INPUT_BRAM_33_DEPTH(C_INPUT_BRAM_33_DEPTH),
        .C_INPUT_BRAM_34_DEPTH(C_INPUT_BRAM_34_DEPTH),
        .C_INPUT_BRAM_35_DEPTH(C_INPUT_BRAM_35_DEPTH),
        .C_INPUT_BRAM_36_DEPTH(C_INPUT_BRAM_36_DEPTH),
        .C_INPUT_BRAM_37_DEPTH(C_INPUT_BRAM_37_DEPTH),
        .C_INPUT_BRAM_38_DEPTH(C_INPUT_BRAM_38_DEPTH),
        .C_INPUT_BRAM_39_DEPTH(C_INPUT_BRAM_39_DEPTH),
        .C_INPUT_BRAM_40_DEPTH(C_INPUT_BRAM_40_DEPTH),
        .C_INPUT_BRAM_41_DEPTH(C_INPUT_BRAM_41_DEPTH),
        .C_INPUT_BRAM_42_DEPTH(C_INPUT_BRAM_42_DEPTH),
        .C_INPUT_BRAM_43_DEPTH(C_INPUT_BRAM_43_DEPTH),
        .C_INPUT_BRAM_44_DEPTH(C_INPUT_BRAM_44_DEPTH),
        .C_INPUT_BRAM_45_DEPTH(C_INPUT_BRAM_45_DEPTH),
        .C_INPUT_BRAM_46_DEPTH(C_INPUT_BRAM_46_DEPTH),
        .C_INPUT_BRAM_47_DEPTH(C_INPUT_BRAM_47_DEPTH),
        .C_INPUT_BRAM_48_DEPTH(C_INPUT_BRAM_48_DEPTH),
        .C_INPUT_BRAM_49_DEPTH(C_INPUT_BRAM_49_DEPTH),
        .C_INPUT_BRAM_50_DEPTH(C_INPUT_BRAM_50_DEPTH),
        .C_INPUT_BRAM_51_DEPTH(C_INPUT_BRAM_51_DEPTH),
        .C_INPUT_BRAM_52_DEPTH(C_INPUT_BRAM_52_DEPTH),
        .C_INPUT_BRAM_53_DEPTH(C_INPUT_BRAM_53_DEPTH),
        .C_INPUT_BRAM_54_DEPTH(C_INPUT_BRAM_54_DEPTH),
        .C_INPUT_BRAM_55_DEPTH(C_INPUT_BRAM_55_DEPTH),
        .C_INPUT_BRAM_56_DEPTH(C_INPUT_BRAM_56_DEPTH),
        .C_INPUT_BRAM_57_DEPTH(C_INPUT_BRAM_57_DEPTH),
        .C_INPUT_BRAM_58_DEPTH(C_INPUT_BRAM_58_DEPTH),
        .C_INPUT_BRAM_59_DEPTH(C_INPUT_BRAM_59_DEPTH),
        .C_INPUT_BRAM_60_DEPTH(C_INPUT_BRAM_60_DEPTH),
        .C_INPUT_BRAM_61_DEPTH(C_INPUT_BRAM_61_DEPTH),
        .C_INPUT_BRAM_62_DEPTH(C_INPUT_BRAM_62_DEPTH),
        .C_INPUT_BRAM_63_DEPTH(C_INPUT_BRAM_63_DEPTH),
        .C_INPUT_BRAM_64_DEPTH(C_INPUT_BRAM_64_DEPTH),
        .C_INPUT_BRAM_65_DEPTH(C_INPUT_BRAM_65_DEPTH),
        .C_INPUT_BRAM_66_DEPTH(C_INPUT_BRAM_66_DEPTH),
        .C_INPUT_BRAM_67_DEPTH(C_INPUT_BRAM_67_DEPTH),
        .C_INPUT_BRAM_68_DEPTH(C_INPUT_BRAM_68_DEPTH),
        .C_INPUT_BRAM_69_DEPTH(C_INPUT_BRAM_69_DEPTH),
        .C_INPUT_BRAM_70_DEPTH(C_INPUT_BRAM_70_DEPTH),
        .C_INPUT_BRAM_71_DEPTH(C_INPUT_BRAM_71_DEPTH),
        .C_INPUT_BRAM_72_DEPTH(C_INPUT_BRAM_72_DEPTH),
        .C_INPUT_BRAM_73_DEPTH(C_INPUT_BRAM_73_DEPTH),
        .C_INPUT_BRAM_74_DEPTH(C_INPUT_BRAM_74_DEPTH),
        .C_INPUT_BRAM_75_DEPTH(C_INPUT_BRAM_75_DEPTH),
        .C_INPUT_BRAM_76_DEPTH(C_INPUT_BRAM_76_DEPTH),
        .C_INPUT_BRAM_77_DEPTH(C_INPUT_BRAM_77_DEPTH),
        .C_INPUT_BRAM_78_DEPTH(C_INPUT_BRAM_78_DEPTH),
        .C_INPUT_BRAM_79_DEPTH(C_INPUT_BRAM_79_DEPTH),
        .C_INPUT_BRAM_80_DEPTH(C_INPUT_BRAM_80_DEPTH),
        .C_INPUT_BRAM_81_DEPTH(C_INPUT_BRAM_81_DEPTH),
        .C_INPUT_BRAM_82_DEPTH(C_INPUT_BRAM_82_DEPTH),
        .C_INPUT_BRAM_83_DEPTH(C_INPUT_BRAM_83_DEPTH),
        .C_INPUT_BRAM_84_DEPTH(C_INPUT_BRAM_84_DEPTH),
        .C_INPUT_BRAM_85_DEPTH(C_INPUT_BRAM_85_DEPTH),
        .C_INPUT_BRAM_86_DEPTH(C_INPUT_BRAM_86_DEPTH),
        .C_INPUT_BRAM_87_DEPTH(C_INPUT_BRAM_87_DEPTH),
        .C_INPUT_BRAM_88_DEPTH(C_INPUT_BRAM_88_DEPTH),
        .C_INPUT_BRAM_89_DEPTH(C_INPUT_BRAM_89_DEPTH),
        .C_INPUT_BRAM_90_DEPTH(C_INPUT_BRAM_90_DEPTH),
        .C_INPUT_BRAM_91_DEPTH(C_INPUT_BRAM_91_DEPTH),
        .C_INPUT_BRAM_92_DEPTH(C_INPUT_BRAM_92_DEPTH),
        .C_INPUT_BRAM_93_DEPTH(C_INPUT_BRAM_93_DEPTH),
        .C_INPUT_BRAM_94_DEPTH(C_INPUT_BRAM_94_DEPTH),
        .C_INPUT_BRAM_95_DEPTH(C_INPUT_BRAM_95_DEPTH),
        .C_INPUT_BRAM_96_DEPTH(C_INPUT_BRAM_96_DEPTH),
        .C_INPUT_BRAM_97_DEPTH(C_INPUT_BRAM_97_DEPTH),
        .C_INPUT_BRAM_98_DEPTH(C_INPUT_BRAM_98_DEPTH),
        .C_INPUT_BRAM_99_DEPTH(C_INPUT_BRAM_99_DEPTH),
        .C_INPUT_BRAM_100_DEPTH(C_INPUT_BRAM_100_DEPTH),
        .C_INPUT_BRAM_101_DEPTH(C_INPUT_BRAM_101_DEPTH),
        .C_INPUT_BRAM_102_DEPTH(C_INPUT_BRAM_102_DEPTH),
        .C_INPUT_BRAM_103_DEPTH(C_INPUT_BRAM_103_DEPTH),
        .C_INPUT_BRAM_104_DEPTH(C_INPUT_BRAM_104_DEPTH),
        .C_INPUT_BRAM_105_DEPTH(C_INPUT_BRAM_105_DEPTH),
        .C_INPUT_BRAM_106_DEPTH(C_INPUT_BRAM_106_DEPTH),
        .C_INPUT_BRAM_107_DEPTH(C_INPUT_BRAM_107_DEPTH),
        .C_INPUT_BRAM_108_DEPTH(C_INPUT_BRAM_108_DEPTH),
        .C_INPUT_BRAM_109_DEPTH(C_INPUT_BRAM_109_DEPTH),
        .C_INPUT_BRAM_110_DEPTH(C_INPUT_BRAM_110_DEPTH),
        .C_INPUT_BRAM_111_DEPTH(C_INPUT_BRAM_111_DEPTH),
        .C_INPUT_BRAM_112_DEPTH(C_INPUT_BRAM_112_DEPTH),
        .C_INPUT_BRAM_113_DEPTH(C_INPUT_BRAM_113_DEPTH),
        .C_INPUT_BRAM_114_DEPTH(C_INPUT_BRAM_114_DEPTH),
        .C_INPUT_BRAM_115_DEPTH(C_INPUT_BRAM_115_DEPTH),
        .C_INPUT_BRAM_116_DEPTH(C_INPUT_BRAM_116_DEPTH),
        .C_INPUT_BRAM_117_DEPTH(C_INPUT_BRAM_117_DEPTH),
        .C_INPUT_BRAM_118_DEPTH(C_INPUT_BRAM_118_DEPTH),
        .C_INPUT_BRAM_119_DEPTH(C_INPUT_BRAM_119_DEPTH),
        .C_INPUT_BRAM_120_DEPTH(C_INPUT_BRAM_120_DEPTH),
        .C_INPUT_BRAM_121_DEPTH(C_INPUT_BRAM_121_DEPTH),
        .C_INPUT_BRAM_122_DEPTH(C_INPUT_BRAM_122_DEPTH),
        .C_INPUT_BRAM_123_DEPTH(C_INPUT_BRAM_123_DEPTH),
        .C_INPUT_BRAM_124_DEPTH(C_INPUT_BRAM_124_DEPTH),
        .C_INPUT_BRAM_125_DEPTH(C_INPUT_BRAM_125_DEPTH),
        .C_INPUT_BRAM_126_DEPTH(C_INPUT_BRAM_126_DEPTH),
        .C_INPUT_BRAM_127_DEPTH(C_INPUT_BRAM_127_DEPTH),
        .C_INPUT_BRAM_0_DMWIDTH(C_INPUT_BRAM_0_DMWIDTH),
        .C_INPUT_BRAM_1_DMWIDTH(C_INPUT_BRAM_1_DMWIDTH),
        .C_INPUT_BRAM_2_DMWIDTH(C_INPUT_BRAM_2_DMWIDTH),
        .C_INPUT_BRAM_3_DMWIDTH(C_INPUT_BRAM_3_DMWIDTH),
        .C_INPUT_BRAM_4_DMWIDTH(C_INPUT_BRAM_4_DMWIDTH),
        .C_INPUT_BRAM_5_DMWIDTH(C_INPUT_BRAM_5_DMWIDTH),
        .C_INPUT_BRAM_6_DMWIDTH(C_INPUT_BRAM_6_DMWIDTH),
        .C_INPUT_BRAM_7_DMWIDTH(C_INPUT_BRAM_7_DMWIDTH),
        .C_INPUT_BRAM_8_DMWIDTH(C_INPUT_BRAM_8_DMWIDTH),
        .C_INPUT_BRAM_9_DMWIDTH(C_INPUT_BRAM_9_DMWIDTH),
        .C_INPUT_BRAM_10_DMWIDTH(C_INPUT_BRAM_10_DMWIDTH),
        .C_INPUT_BRAM_11_DMWIDTH(C_INPUT_BRAM_11_DMWIDTH),
        .C_INPUT_BRAM_12_DMWIDTH(C_INPUT_BRAM_12_DMWIDTH),
        .C_INPUT_BRAM_13_DMWIDTH(C_INPUT_BRAM_13_DMWIDTH),
        .C_INPUT_BRAM_14_DMWIDTH(C_INPUT_BRAM_14_DMWIDTH),
        .C_INPUT_BRAM_15_DMWIDTH(C_INPUT_BRAM_15_DMWIDTH),
        .C_INPUT_BRAM_16_DMWIDTH(C_INPUT_BRAM_16_DMWIDTH),
        .C_INPUT_BRAM_17_DMWIDTH(C_INPUT_BRAM_17_DMWIDTH),
        .C_INPUT_BRAM_18_DMWIDTH(C_INPUT_BRAM_18_DMWIDTH),
        .C_INPUT_BRAM_19_DMWIDTH(C_INPUT_BRAM_19_DMWIDTH),
        .C_INPUT_BRAM_20_DMWIDTH(C_INPUT_BRAM_20_DMWIDTH),
        .C_INPUT_BRAM_21_DMWIDTH(C_INPUT_BRAM_21_DMWIDTH),
        .C_INPUT_BRAM_22_DMWIDTH(C_INPUT_BRAM_22_DMWIDTH),
        .C_INPUT_BRAM_23_DMWIDTH(C_INPUT_BRAM_23_DMWIDTH),
        .C_INPUT_BRAM_24_DMWIDTH(C_INPUT_BRAM_24_DMWIDTH),
        .C_INPUT_BRAM_25_DMWIDTH(C_INPUT_BRAM_25_DMWIDTH),
        .C_INPUT_BRAM_26_DMWIDTH(C_INPUT_BRAM_26_DMWIDTH),
        .C_INPUT_BRAM_27_DMWIDTH(C_INPUT_BRAM_27_DMWIDTH),
        .C_INPUT_BRAM_28_DMWIDTH(C_INPUT_BRAM_28_DMWIDTH),
        .C_INPUT_BRAM_29_DMWIDTH(C_INPUT_BRAM_29_DMWIDTH),
        .C_INPUT_BRAM_30_DMWIDTH(C_INPUT_BRAM_30_DMWIDTH),
        .C_INPUT_BRAM_31_DMWIDTH(C_INPUT_BRAM_31_DMWIDTH),
        .C_INPUT_BRAM_32_DMWIDTH(C_INPUT_BRAM_32_DMWIDTH),
        .C_INPUT_BRAM_33_DMWIDTH(C_INPUT_BRAM_33_DMWIDTH),
        .C_INPUT_BRAM_34_DMWIDTH(C_INPUT_BRAM_34_DMWIDTH),
        .C_INPUT_BRAM_35_DMWIDTH(C_INPUT_BRAM_35_DMWIDTH),
        .C_INPUT_BRAM_36_DMWIDTH(C_INPUT_BRAM_36_DMWIDTH),
        .C_INPUT_BRAM_37_DMWIDTH(C_INPUT_BRAM_37_DMWIDTH),
        .C_INPUT_BRAM_38_DMWIDTH(C_INPUT_BRAM_38_DMWIDTH),
        .C_INPUT_BRAM_39_DMWIDTH(C_INPUT_BRAM_39_DMWIDTH),
        .C_INPUT_BRAM_40_DMWIDTH(C_INPUT_BRAM_40_DMWIDTH),
        .C_INPUT_BRAM_41_DMWIDTH(C_INPUT_BRAM_41_DMWIDTH),
        .C_INPUT_BRAM_42_DMWIDTH(C_INPUT_BRAM_42_DMWIDTH),
        .C_INPUT_BRAM_43_DMWIDTH(C_INPUT_BRAM_43_DMWIDTH),
        .C_INPUT_BRAM_44_DMWIDTH(C_INPUT_BRAM_44_DMWIDTH),
        .C_INPUT_BRAM_45_DMWIDTH(C_INPUT_BRAM_45_DMWIDTH),
        .C_INPUT_BRAM_46_DMWIDTH(C_INPUT_BRAM_46_DMWIDTH),
        .C_INPUT_BRAM_47_DMWIDTH(C_INPUT_BRAM_47_DMWIDTH),
        .C_INPUT_BRAM_48_DMWIDTH(C_INPUT_BRAM_48_DMWIDTH),
        .C_INPUT_BRAM_49_DMWIDTH(C_INPUT_BRAM_49_DMWIDTH),
        .C_INPUT_BRAM_50_DMWIDTH(C_INPUT_BRAM_50_DMWIDTH),
        .C_INPUT_BRAM_51_DMWIDTH(C_INPUT_BRAM_51_DMWIDTH),
        .C_INPUT_BRAM_52_DMWIDTH(C_INPUT_BRAM_52_DMWIDTH),
        .C_INPUT_BRAM_53_DMWIDTH(C_INPUT_BRAM_53_DMWIDTH),
        .C_INPUT_BRAM_54_DMWIDTH(C_INPUT_BRAM_54_DMWIDTH),
        .C_INPUT_BRAM_55_DMWIDTH(C_INPUT_BRAM_55_DMWIDTH),
        .C_INPUT_BRAM_56_DMWIDTH(C_INPUT_BRAM_56_DMWIDTH),
        .C_INPUT_BRAM_57_DMWIDTH(C_INPUT_BRAM_57_DMWIDTH),
        .C_INPUT_BRAM_58_DMWIDTH(C_INPUT_BRAM_58_DMWIDTH),
        .C_INPUT_BRAM_59_DMWIDTH(C_INPUT_BRAM_59_DMWIDTH),
        .C_INPUT_BRAM_60_DMWIDTH(C_INPUT_BRAM_60_DMWIDTH),
        .C_INPUT_BRAM_61_DMWIDTH(C_INPUT_BRAM_61_DMWIDTH),
        .C_INPUT_BRAM_62_DMWIDTH(C_INPUT_BRAM_62_DMWIDTH),
        .C_INPUT_BRAM_63_DMWIDTH(C_INPUT_BRAM_63_DMWIDTH),
        .C_INPUT_BRAM_64_DMWIDTH(C_INPUT_BRAM_64_DMWIDTH),
        .C_INPUT_BRAM_65_DMWIDTH(C_INPUT_BRAM_65_DMWIDTH),
        .C_INPUT_BRAM_66_DMWIDTH(C_INPUT_BRAM_66_DMWIDTH),
        .C_INPUT_BRAM_67_DMWIDTH(C_INPUT_BRAM_67_DMWIDTH),
        .C_INPUT_BRAM_68_DMWIDTH(C_INPUT_BRAM_68_DMWIDTH),
        .C_INPUT_BRAM_69_DMWIDTH(C_INPUT_BRAM_69_DMWIDTH),
        .C_INPUT_BRAM_70_DMWIDTH(C_INPUT_BRAM_70_DMWIDTH),
        .C_INPUT_BRAM_71_DMWIDTH(C_INPUT_BRAM_71_DMWIDTH),
        .C_INPUT_BRAM_72_DMWIDTH(C_INPUT_BRAM_72_DMWIDTH),
        .C_INPUT_BRAM_73_DMWIDTH(C_INPUT_BRAM_73_DMWIDTH),
        .C_INPUT_BRAM_74_DMWIDTH(C_INPUT_BRAM_74_DMWIDTH),
        .C_INPUT_BRAM_75_DMWIDTH(C_INPUT_BRAM_75_DMWIDTH),
        .C_INPUT_BRAM_76_DMWIDTH(C_INPUT_BRAM_76_DMWIDTH),
        .C_INPUT_BRAM_77_DMWIDTH(C_INPUT_BRAM_77_DMWIDTH),
        .C_INPUT_BRAM_78_DMWIDTH(C_INPUT_BRAM_78_DMWIDTH),
        .C_INPUT_BRAM_79_DMWIDTH(C_INPUT_BRAM_79_DMWIDTH),
        .C_INPUT_BRAM_80_DMWIDTH(C_INPUT_BRAM_80_DMWIDTH),
        .C_INPUT_BRAM_81_DMWIDTH(C_INPUT_BRAM_81_DMWIDTH),
        .C_INPUT_BRAM_82_DMWIDTH(C_INPUT_BRAM_82_DMWIDTH),
        .C_INPUT_BRAM_83_DMWIDTH(C_INPUT_BRAM_83_DMWIDTH),
        .C_INPUT_BRAM_84_DMWIDTH(C_INPUT_BRAM_84_DMWIDTH),
        .C_INPUT_BRAM_85_DMWIDTH(C_INPUT_BRAM_85_DMWIDTH),
        .C_INPUT_BRAM_86_DMWIDTH(C_INPUT_BRAM_86_DMWIDTH),
        .C_INPUT_BRAM_87_DMWIDTH(C_INPUT_BRAM_87_DMWIDTH),
        .C_INPUT_BRAM_88_DMWIDTH(C_INPUT_BRAM_88_DMWIDTH),
        .C_INPUT_BRAM_89_DMWIDTH(C_INPUT_BRAM_89_DMWIDTH),
        .C_INPUT_BRAM_90_DMWIDTH(C_INPUT_BRAM_90_DMWIDTH),
        .C_INPUT_BRAM_91_DMWIDTH(C_INPUT_BRAM_91_DMWIDTH),
        .C_INPUT_BRAM_92_DMWIDTH(C_INPUT_BRAM_92_DMWIDTH),
        .C_INPUT_BRAM_93_DMWIDTH(C_INPUT_BRAM_93_DMWIDTH),
        .C_INPUT_BRAM_94_DMWIDTH(C_INPUT_BRAM_94_DMWIDTH),
        .C_INPUT_BRAM_95_DMWIDTH(C_INPUT_BRAM_95_DMWIDTH),
        .C_INPUT_BRAM_96_DMWIDTH(C_INPUT_BRAM_96_DMWIDTH),
        .C_INPUT_BRAM_97_DMWIDTH(C_INPUT_BRAM_97_DMWIDTH),
        .C_INPUT_BRAM_98_DMWIDTH(C_INPUT_BRAM_98_DMWIDTH),
        .C_INPUT_BRAM_99_DMWIDTH(C_INPUT_BRAM_99_DMWIDTH),
        .C_INPUT_BRAM_100_DMWIDTH(C_INPUT_BRAM_100_DMWIDTH),
        .C_INPUT_BRAM_101_DMWIDTH(C_INPUT_BRAM_101_DMWIDTH),
        .C_INPUT_BRAM_102_DMWIDTH(C_INPUT_BRAM_102_DMWIDTH),
        .C_INPUT_BRAM_103_DMWIDTH(C_INPUT_BRAM_103_DMWIDTH),
        .C_INPUT_BRAM_104_DMWIDTH(C_INPUT_BRAM_104_DMWIDTH),
        .C_INPUT_BRAM_105_DMWIDTH(C_INPUT_BRAM_105_DMWIDTH),
        .C_INPUT_BRAM_106_DMWIDTH(C_INPUT_BRAM_106_DMWIDTH),
        .C_INPUT_BRAM_107_DMWIDTH(C_INPUT_BRAM_107_DMWIDTH),
        .C_INPUT_BRAM_108_DMWIDTH(C_INPUT_BRAM_108_DMWIDTH),
        .C_INPUT_BRAM_109_DMWIDTH(C_INPUT_BRAM_109_DMWIDTH),
        .C_INPUT_BRAM_110_DMWIDTH(C_INPUT_BRAM_110_DMWIDTH),
        .C_INPUT_BRAM_111_DMWIDTH(C_INPUT_BRAM_111_DMWIDTH),
        .C_INPUT_BRAM_112_DMWIDTH(C_INPUT_BRAM_112_DMWIDTH),
        .C_INPUT_BRAM_113_DMWIDTH(C_INPUT_BRAM_113_DMWIDTH),
        .C_INPUT_BRAM_114_DMWIDTH(C_INPUT_BRAM_114_DMWIDTH),
        .C_INPUT_BRAM_115_DMWIDTH(C_INPUT_BRAM_115_DMWIDTH),
        .C_INPUT_BRAM_116_DMWIDTH(C_INPUT_BRAM_116_DMWIDTH),
        .C_INPUT_BRAM_117_DMWIDTH(C_INPUT_BRAM_117_DMWIDTH),
        .C_INPUT_BRAM_118_DMWIDTH(C_INPUT_BRAM_118_DMWIDTH),
        .C_INPUT_BRAM_119_DMWIDTH(C_INPUT_BRAM_119_DMWIDTH),
        .C_INPUT_BRAM_120_DMWIDTH(C_INPUT_BRAM_120_DMWIDTH),
        .C_INPUT_BRAM_121_DMWIDTH(C_INPUT_BRAM_121_DMWIDTH),
        .C_INPUT_BRAM_122_DMWIDTH(C_INPUT_BRAM_122_DMWIDTH),
        .C_INPUT_BRAM_123_DMWIDTH(C_INPUT_BRAM_123_DMWIDTH),
        .C_INPUT_BRAM_124_DMWIDTH(C_INPUT_BRAM_124_DMWIDTH),
        .C_INPUT_BRAM_125_DMWIDTH(C_INPUT_BRAM_125_DMWIDTH),
        .C_INPUT_BRAM_126_DMWIDTH(C_INPUT_BRAM_126_DMWIDTH),
        .C_INPUT_BRAM_127_DMWIDTH(C_INPUT_BRAM_127_DMWIDTH),
        .C_OUTPUT_BRAM_0_DMWIDTH(C_INOUT_BRAM_0_DMWIDTH),
        .C_OUTPUT_BRAM_1_DMWIDTH(C_INOUT_BRAM_1_DMWIDTH),
        .C_OUTPUT_BRAM_2_DMWIDTH(C_INOUT_BRAM_2_DMWIDTH),
        .C_OUTPUT_BRAM_3_DMWIDTH(C_INOUT_BRAM_3_DMWIDTH),
        .C_OUTPUT_BRAM_4_DMWIDTH(C_INOUT_BRAM_4_DMWIDTH),
        .C_OUTPUT_BRAM_5_DMWIDTH(C_INOUT_BRAM_5_DMWIDTH),
        .C_OUTPUT_BRAM_6_DMWIDTH(C_INOUT_BRAM_6_DMWIDTH),
        .C_OUTPUT_BRAM_7_DMWIDTH(C_INOUT_BRAM_7_DMWIDTH),
        .C_OUTPUT_BRAM_8_DMWIDTH(C_INOUT_BRAM_8_DMWIDTH),
        .C_OUTPUT_BRAM_9_DMWIDTH(C_INOUT_BRAM_9_DMWIDTH),
        .C_OUTPUT_BRAM_10_DMWIDTH(C_INOUT_BRAM_10_DMWIDTH),
        .C_OUTPUT_BRAM_11_DMWIDTH(C_INOUT_BRAM_11_DMWIDTH),
        .C_OUTPUT_BRAM_12_DMWIDTH(C_INOUT_BRAM_12_DMWIDTH),
        .C_OUTPUT_BRAM_13_DMWIDTH(C_INOUT_BRAM_13_DMWIDTH),
        .C_OUTPUT_BRAM_14_DMWIDTH(C_INOUT_BRAM_14_DMWIDTH),
        .C_OUTPUT_BRAM_15_DMWIDTH(C_INOUT_BRAM_15_DMWIDTH),
        .C_OUTPUT_BRAM_16_DMWIDTH(C_INOUT_BRAM_16_DMWIDTH),
        .C_OUTPUT_BRAM_17_DMWIDTH(C_INOUT_BRAM_17_DMWIDTH),
        .C_OUTPUT_BRAM_18_DMWIDTH(C_INOUT_BRAM_18_DMWIDTH),
        .C_OUTPUT_BRAM_19_DMWIDTH(C_INOUT_BRAM_19_DMWIDTH),
        .C_OUTPUT_BRAM_20_DMWIDTH(C_INOUT_BRAM_20_DMWIDTH),
        .C_OUTPUT_BRAM_21_DMWIDTH(C_INOUT_BRAM_21_DMWIDTH),
        .C_OUTPUT_BRAM_22_DMWIDTH(C_INOUT_BRAM_22_DMWIDTH),
        .C_OUTPUT_BRAM_23_DMWIDTH(C_INOUT_BRAM_23_DMWIDTH),
        .C_OUTPUT_BRAM_24_DMWIDTH(C_INOUT_BRAM_24_DMWIDTH),
        .C_OUTPUT_BRAM_25_DMWIDTH(C_INOUT_BRAM_25_DMWIDTH),
        .C_OUTPUT_BRAM_26_DMWIDTH(C_INOUT_BRAM_26_DMWIDTH),
        .C_OUTPUT_BRAM_27_DMWIDTH(C_INOUT_BRAM_27_DMWIDTH),
        .C_OUTPUT_BRAM_28_DMWIDTH(C_INOUT_BRAM_28_DMWIDTH),
        .C_OUTPUT_BRAM_29_DMWIDTH(C_INOUT_BRAM_29_DMWIDTH),
        .C_OUTPUT_BRAM_30_DMWIDTH(C_INOUT_BRAM_30_DMWIDTH),
        .C_OUTPUT_BRAM_31_DMWIDTH(C_INOUT_BRAM_31_DMWIDTH),
        .C_OUTPUT_BRAM_32_DMWIDTH(C_INOUT_BRAM_32_DMWIDTH),
        .C_OUTPUT_BRAM_33_DMWIDTH(C_INOUT_BRAM_33_DMWIDTH),
        .C_OUTPUT_BRAM_34_DMWIDTH(C_INOUT_BRAM_34_DMWIDTH),
        .C_OUTPUT_BRAM_35_DMWIDTH(C_INOUT_BRAM_35_DMWIDTH),
        .C_OUTPUT_BRAM_36_DMWIDTH(C_INOUT_BRAM_36_DMWIDTH),
        .C_OUTPUT_BRAM_37_DMWIDTH(C_INOUT_BRAM_37_DMWIDTH),
        .C_OUTPUT_BRAM_38_DMWIDTH(C_INOUT_BRAM_38_DMWIDTH),
        .C_OUTPUT_BRAM_39_DMWIDTH(C_INOUT_BRAM_39_DMWIDTH),
        .C_OUTPUT_BRAM_40_DMWIDTH(C_INOUT_BRAM_40_DMWIDTH),
        .C_OUTPUT_BRAM_41_DMWIDTH(C_INOUT_BRAM_41_DMWIDTH),
        .C_OUTPUT_BRAM_42_DMWIDTH(C_INOUT_BRAM_42_DMWIDTH),
        .C_OUTPUT_BRAM_43_DMWIDTH(C_INOUT_BRAM_43_DMWIDTH),
        .C_OUTPUT_BRAM_44_DMWIDTH(C_INOUT_BRAM_44_DMWIDTH),
        .C_OUTPUT_BRAM_45_DMWIDTH(C_INOUT_BRAM_45_DMWIDTH),
        .C_OUTPUT_BRAM_46_DMWIDTH(C_INOUT_BRAM_46_DMWIDTH),
        .C_OUTPUT_BRAM_47_DMWIDTH(C_INOUT_BRAM_47_DMWIDTH),
        .C_OUTPUT_BRAM_48_DMWIDTH(C_INOUT_BRAM_48_DMWIDTH),
        .C_OUTPUT_BRAM_49_DMWIDTH(C_INOUT_BRAM_49_DMWIDTH),
        .C_OUTPUT_BRAM_50_DMWIDTH(C_INOUT_BRAM_50_DMWIDTH),
        .C_OUTPUT_BRAM_51_DMWIDTH(C_INOUT_BRAM_51_DMWIDTH),
        .C_OUTPUT_BRAM_52_DMWIDTH(C_INOUT_BRAM_52_DMWIDTH),
        .C_OUTPUT_BRAM_53_DMWIDTH(C_INOUT_BRAM_53_DMWIDTH),
        .C_OUTPUT_BRAM_54_DMWIDTH(C_INOUT_BRAM_54_DMWIDTH),
        .C_OUTPUT_BRAM_55_DMWIDTH(C_INOUT_BRAM_55_DMWIDTH),
        .C_OUTPUT_BRAM_56_DMWIDTH(C_INOUT_BRAM_56_DMWIDTH),
        .C_OUTPUT_BRAM_57_DMWIDTH(C_INOUT_BRAM_57_DMWIDTH),
        .C_OUTPUT_BRAM_58_DMWIDTH(C_INOUT_BRAM_58_DMWIDTH),
        .C_OUTPUT_BRAM_59_DMWIDTH(C_INOUT_BRAM_59_DMWIDTH),
        .C_OUTPUT_BRAM_60_DMWIDTH(C_INOUT_BRAM_60_DMWIDTH),
        .C_OUTPUT_BRAM_61_DMWIDTH(C_INOUT_BRAM_61_DMWIDTH),
        .C_OUTPUT_BRAM_62_DMWIDTH(C_INOUT_BRAM_62_DMWIDTH),
        .C_OUTPUT_BRAM_63_DMWIDTH(C_INOUT_BRAM_63_DMWIDTH),
        .C_OUTPUT_BRAM_64_DMWIDTH(C_INOUT_BRAM_64_DMWIDTH),
        .C_OUTPUT_BRAM_65_DMWIDTH(C_INOUT_BRAM_65_DMWIDTH),
        .C_OUTPUT_BRAM_66_DMWIDTH(C_INOUT_BRAM_66_DMWIDTH),
        .C_OUTPUT_BRAM_67_DMWIDTH(C_INOUT_BRAM_67_DMWIDTH),
        .C_OUTPUT_BRAM_68_DMWIDTH(C_INOUT_BRAM_68_DMWIDTH),
        .C_OUTPUT_BRAM_69_DMWIDTH(C_INOUT_BRAM_69_DMWIDTH),
        .C_OUTPUT_BRAM_70_DMWIDTH(C_INOUT_BRAM_70_DMWIDTH),
        .C_OUTPUT_BRAM_71_DMWIDTH(C_INOUT_BRAM_71_DMWIDTH),
        .C_OUTPUT_BRAM_72_DMWIDTH(C_INOUT_BRAM_72_DMWIDTH),
        .C_OUTPUT_BRAM_73_DMWIDTH(C_INOUT_BRAM_73_DMWIDTH),
        .C_OUTPUT_BRAM_74_DMWIDTH(C_INOUT_BRAM_74_DMWIDTH),
        .C_OUTPUT_BRAM_75_DMWIDTH(C_INOUT_BRAM_75_DMWIDTH),
        .C_OUTPUT_BRAM_76_DMWIDTH(C_INOUT_BRAM_76_DMWIDTH),
        .C_OUTPUT_BRAM_77_DMWIDTH(C_INOUT_BRAM_77_DMWIDTH),
        .C_OUTPUT_BRAM_78_DMWIDTH(C_INOUT_BRAM_78_DMWIDTH),
        .C_OUTPUT_BRAM_79_DMWIDTH(C_INOUT_BRAM_79_DMWIDTH),
        .C_OUTPUT_BRAM_80_DMWIDTH(C_INOUT_BRAM_80_DMWIDTH),
        .C_OUTPUT_BRAM_81_DMWIDTH(C_INOUT_BRAM_81_DMWIDTH),
        .C_OUTPUT_BRAM_82_DMWIDTH(C_INOUT_BRAM_82_DMWIDTH),
        .C_OUTPUT_BRAM_83_DMWIDTH(C_INOUT_BRAM_83_DMWIDTH),
        .C_OUTPUT_BRAM_84_DMWIDTH(C_INOUT_BRAM_84_DMWIDTH),
        .C_OUTPUT_BRAM_85_DMWIDTH(C_INOUT_BRAM_85_DMWIDTH),
        .C_OUTPUT_BRAM_86_DMWIDTH(C_INOUT_BRAM_86_DMWIDTH),
        .C_OUTPUT_BRAM_87_DMWIDTH(C_INOUT_BRAM_87_DMWIDTH),
        .C_OUTPUT_BRAM_88_DMWIDTH(C_INOUT_BRAM_88_DMWIDTH),
        .C_OUTPUT_BRAM_89_DMWIDTH(C_INOUT_BRAM_89_DMWIDTH),
        .C_OUTPUT_BRAM_90_DMWIDTH(C_INOUT_BRAM_90_DMWIDTH),
        .C_OUTPUT_BRAM_91_DMWIDTH(C_INOUT_BRAM_91_DMWIDTH),
        .C_OUTPUT_BRAM_92_DMWIDTH(C_INOUT_BRAM_92_DMWIDTH),
        .C_OUTPUT_BRAM_93_DMWIDTH(C_INOUT_BRAM_93_DMWIDTH),
        .C_OUTPUT_BRAM_94_DMWIDTH(C_INOUT_BRAM_94_DMWIDTH),
        .C_OUTPUT_BRAM_95_DMWIDTH(C_INOUT_BRAM_95_DMWIDTH),
        .C_OUTPUT_BRAM_96_DMWIDTH(C_INOUT_BRAM_96_DMWIDTH),
        .C_OUTPUT_BRAM_97_DMWIDTH(C_INOUT_BRAM_97_DMWIDTH),
        .C_OUTPUT_BRAM_98_DMWIDTH(C_INOUT_BRAM_98_DMWIDTH),
        .C_OUTPUT_BRAM_99_DMWIDTH(C_INOUT_BRAM_99_DMWIDTH),
        .C_OUTPUT_BRAM_100_DMWIDTH(C_INOUT_BRAM_100_DMWIDTH),
        .C_OUTPUT_BRAM_101_DMWIDTH(C_INOUT_BRAM_101_DMWIDTH),
        .C_OUTPUT_BRAM_102_DMWIDTH(C_INOUT_BRAM_102_DMWIDTH),
        .C_OUTPUT_BRAM_103_DMWIDTH(C_INOUT_BRAM_103_DMWIDTH),
        .C_OUTPUT_BRAM_104_DMWIDTH(C_INOUT_BRAM_104_DMWIDTH),
        .C_OUTPUT_BRAM_105_DMWIDTH(C_INOUT_BRAM_105_DMWIDTH),
        .C_OUTPUT_BRAM_106_DMWIDTH(C_INOUT_BRAM_106_DMWIDTH),
        .C_OUTPUT_BRAM_107_DMWIDTH(C_INOUT_BRAM_107_DMWIDTH),
        .C_OUTPUT_BRAM_108_DMWIDTH(C_INOUT_BRAM_108_DMWIDTH),
        .C_OUTPUT_BRAM_109_DMWIDTH(C_INOUT_BRAM_109_DMWIDTH),
        .C_OUTPUT_BRAM_110_DMWIDTH(C_INOUT_BRAM_110_DMWIDTH),
        .C_OUTPUT_BRAM_111_DMWIDTH(C_INOUT_BRAM_111_DMWIDTH),
        .C_OUTPUT_BRAM_112_DMWIDTH(C_INOUT_BRAM_112_DMWIDTH),
        .C_OUTPUT_BRAM_113_DMWIDTH(C_INOUT_BRAM_113_DMWIDTH),
        .C_OUTPUT_BRAM_114_DMWIDTH(C_INOUT_BRAM_114_DMWIDTH),
        .C_OUTPUT_BRAM_115_DMWIDTH(C_INOUT_BRAM_115_DMWIDTH),
        .C_OUTPUT_BRAM_116_DMWIDTH(C_INOUT_BRAM_116_DMWIDTH),
        .C_OUTPUT_BRAM_117_DMWIDTH(C_INOUT_BRAM_117_DMWIDTH),
        .C_OUTPUT_BRAM_118_DMWIDTH(C_INOUT_BRAM_118_DMWIDTH),
        .C_OUTPUT_BRAM_119_DMWIDTH(C_INOUT_BRAM_119_DMWIDTH),
        .C_OUTPUT_BRAM_120_DMWIDTH(C_INOUT_BRAM_120_DMWIDTH),
        .C_OUTPUT_BRAM_121_DMWIDTH(C_INOUT_BRAM_121_DMWIDTH),
        .C_OUTPUT_BRAM_122_DMWIDTH(C_INOUT_BRAM_122_DMWIDTH),
        .C_OUTPUT_BRAM_123_DMWIDTH(C_INOUT_BRAM_123_DMWIDTH),
        .C_OUTPUT_BRAM_124_DMWIDTH(C_INOUT_BRAM_124_DMWIDTH),
        .C_OUTPUT_BRAM_125_DMWIDTH(C_INOUT_BRAM_125_DMWIDTH),
        .C_OUTPUT_BRAM_126_DMWIDTH(C_INOUT_BRAM_126_DMWIDTH),
        .C_OUTPUT_BRAM_127_DMWIDTH(C_INOUT_BRAM_127_DMWIDTH),
        .C_BRAM_0_IS_INOUT(C_BRAM_0_IS_INOUT),
        .C_BRAM_1_IS_INOUT(C_BRAM_1_IS_INOUT),
        .C_BRAM_2_IS_INOUT(C_BRAM_2_IS_INOUT),
        .C_BRAM_3_IS_INOUT(C_BRAM_3_IS_INOUT),
        .C_BRAM_4_IS_INOUT(C_BRAM_4_IS_INOUT),
        .C_BRAM_5_IS_INOUT(C_BRAM_5_IS_INOUT),
        .C_BRAM_6_IS_INOUT(C_BRAM_6_IS_INOUT),
        .C_BRAM_7_IS_INOUT(C_BRAM_7_IS_INOUT),
        .C_BRAM_8_IS_INOUT(C_BRAM_8_IS_INOUT),
        .C_BRAM_9_IS_INOUT(C_BRAM_9_IS_INOUT),
        .C_BRAM_10_IS_INOUT(C_BRAM_10_IS_INOUT),
        .C_BRAM_11_IS_INOUT(C_BRAM_11_IS_INOUT),
        .C_BRAM_12_IS_INOUT(C_BRAM_12_IS_INOUT),
        .C_BRAM_13_IS_INOUT(C_BRAM_13_IS_INOUT),
        .C_BRAM_14_IS_INOUT(C_BRAM_14_IS_INOUT),
        .C_BRAM_15_IS_INOUT(C_BRAM_15_IS_INOUT),
        .C_BRAM_16_IS_INOUT(C_BRAM_16_IS_INOUT),
        .C_BRAM_17_IS_INOUT(C_BRAM_17_IS_INOUT),
        .C_BRAM_18_IS_INOUT(C_BRAM_18_IS_INOUT),
        .C_BRAM_19_IS_INOUT(C_BRAM_19_IS_INOUT),
        .C_BRAM_20_IS_INOUT(C_BRAM_20_IS_INOUT),
        .C_BRAM_21_IS_INOUT(C_BRAM_21_IS_INOUT),
        .C_BRAM_22_IS_INOUT(C_BRAM_22_IS_INOUT),
        .C_BRAM_23_IS_INOUT(C_BRAM_23_IS_INOUT),
        .C_BRAM_24_IS_INOUT(C_BRAM_24_IS_INOUT),
        .C_BRAM_25_IS_INOUT(C_BRAM_25_IS_INOUT),
        .C_BRAM_26_IS_INOUT(C_BRAM_26_IS_INOUT),
        .C_BRAM_27_IS_INOUT(C_BRAM_27_IS_INOUT),
        .C_BRAM_28_IS_INOUT(C_BRAM_28_IS_INOUT),
        .C_BRAM_29_IS_INOUT(C_BRAM_29_IS_INOUT),
        .C_BRAM_30_IS_INOUT(C_BRAM_30_IS_INOUT),
        .C_BRAM_31_IS_INOUT(C_BRAM_31_IS_INOUT),
        .C_BRAM_32_IS_INOUT(C_BRAM_32_IS_INOUT),
        .C_BRAM_33_IS_INOUT(C_BRAM_33_IS_INOUT),
        .C_BRAM_34_IS_INOUT(C_BRAM_34_IS_INOUT),
        .C_BRAM_35_IS_INOUT(C_BRAM_35_IS_INOUT),
        .C_BRAM_36_IS_INOUT(C_BRAM_36_IS_INOUT),
        .C_BRAM_37_IS_INOUT(C_BRAM_37_IS_INOUT),
        .C_BRAM_38_IS_INOUT(C_BRAM_38_IS_INOUT),
        .C_BRAM_39_IS_INOUT(C_BRAM_39_IS_INOUT),
        .C_BRAM_40_IS_INOUT(C_BRAM_40_IS_INOUT),
        .C_BRAM_41_IS_INOUT(C_BRAM_41_IS_INOUT),
        .C_BRAM_42_IS_INOUT(C_BRAM_42_IS_INOUT),
        .C_BRAM_43_IS_INOUT(C_BRAM_43_IS_INOUT),
        .C_BRAM_44_IS_INOUT(C_BRAM_44_IS_INOUT),
        .C_BRAM_45_IS_INOUT(C_BRAM_45_IS_INOUT),
        .C_BRAM_46_IS_INOUT(C_BRAM_46_IS_INOUT),
        .C_BRAM_47_IS_INOUT(C_BRAM_47_IS_INOUT),
        .C_BRAM_48_IS_INOUT(C_BRAM_48_IS_INOUT),
        .C_BRAM_49_IS_INOUT(C_BRAM_49_IS_INOUT),
        .C_BRAM_50_IS_INOUT(C_BRAM_50_IS_INOUT),
        .C_BRAM_51_IS_INOUT(C_BRAM_51_IS_INOUT),
        .C_BRAM_52_IS_INOUT(C_BRAM_52_IS_INOUT),
        .C_BRAM_53_IS_INOUT(C_BRAM_53_IS_INOUT),
        .C_BRAM_54_IS_INOUT(C_BRAM_54_IS_INOUT),
        .C_BRAM_55_IS_INOUT(C_BRAM_55_IS_INOUT),
        .C_BRAM_56_IS_INOUT(C_BRAM_56_IS_INOUT),
        .C_BRAM_57_IS_INOUT(C_BRAM_57_IS_INOUT),
        .C_BRAM_58_IS_INOUT(C_BRAM_58_IS_INOUT),
        .C_BRAM_59_IS_INOUT(C_BRAM_59_IS_INOUT),
        .C_BRAM_60_IS_INOUT(C_BRAM_60_IS_INOUT),
        .C_BRAM_61_IS_INOUT(C_BRAM_61_IS_INOUT),
        .C_BRAM_62_IS_INOUT(C_BRAM_62_IS_INOUT),
        .C_BRAM_63_IS_INOUT(C_BRAM_63_IS_INOUT),
        .C_BRAM_64_IS_INOUT(C_BRAM_64_IS_INOUT),
        .C_BRAM_65_IS_INOUT(C_BRAM_65_IS_INOUT),
        .C_BRAM_66_IS_INOUT(C_BRAM_66_IS_INOUT),
        .C_BRAM_67_IS_INOUT(C_BRAM_67_IS_INOUT),
        .C_BRAM_68_IS_INOUT(C_BRAM_68_IS_INOUT),
        .C_BRAM_69_IS_INOUT(C_BRAM_69_IS_INOUT),
        .C_BRAM_70_IS_INOUT(C_BRAM_70_IS_INOUT),
        .C_BRAM_71_IS_INOUT(C_BRAM_71_IS_INOUT),
        .C_BRAM_72_IS_INOUT(C_BRAM_72_IS_INOUT),
        .C_BRAM_73_IS_INOUT(C_BRAM_73_IS_INOUT),
        .C_BRAM_74_IS_INOUT(C_BRAM_74_IS_INOUT),
        .C_BRAM_75_IS_INOUT(C_BRAM_75_IS_INOUT),
        .C_BRAM_76_IS_INOUT(C_BRAM_76_IS_INOUT),
        .C_BRAM_77_IS_INOUT(C_BRAM_77_IS_INOUT),
        .C_BRAM_78_IS_INOUT(C_BRAM_78_IS_INOUT),
        .C_BRAM_79_IS_INOUT(C_BRAM_79_IS_INOUT),
        .C_BRAM_80_IS_INOUT(C_BRAM_80_IS_INOUT),
        .C_BRAM_81_IS_INOUT(C_BRAM_81_IS_INOUT),
        .C_BRAM_82_IS_INOUT(C_BRAM_82_IS_INOUT),
        .C_BRAM_83_IS_INOUT(C_BRAM_83_IS_INOUT),
        .C_BRAM_84_IS_INOUT(C_BRAM_84_IS_INOUT),
        .C_BRAM_85_IS_INOUT(C_BRAM_85_IS_INOUT),
        .C_BRAM_86_IS_INOUT(C_BRAM_86_IS_INOUT),
        .C_BRAM_87_IS_INOUT(C_BRAM_87_IS_INOUT),
        .C_BRAM_88_IS_INOUT(C_BRAM_88_IS_INOUT),
        .C_BRAM_89_IS_INOUT(C_BRAM_89_IS_INOUT),
        .C_BRAM_90_IS_INOUT(C_BRAM_90_IS_INOUT),
        .C_BRAM_91_IS_INOUT(C_BRAM_91_IS_INOUT),
        .C_BRAM_92_IS_INOUT(C_BRAM_92_IS_INOUT),
        .C_BRAM_93_IS_INOUT(C_BRAM_93_IS_INOUT),
        .C_BRAM_94_IS_INOUT(C_BRAM_94_IS_INOUT),
        .C_BRAM_95_IS_INOUT(C_BRAM_95_IS_INOUT),
        .C_BRAM_96_IS_INOUT(C_BRAM_96_IS_INOUT),
        .C_BRAM_97_IS_INOUT(C_BRAM_97_IS_INOUT),
        .C_BRAM_98_IS_INOUT(C_BRAM_98_IS_INOUT),
        .C_BRAM_99_IS_INOUT(C_BRAM_99_IS_INOUT),
        .C_BRAM_100_IS_INOUT(C_BRAM_100_IS_INOUT),
        .C_BRAM_101_IS_INOUT(C_BRAM_101_IS_INOUT),
        .C_BRAM_102_IS_INOUT(C_BRAM_102_IS_INOUT),
        .C_BRAM_103_IS_INOUT(C_BRAM_103_IS_INOUT),
        .C_BRAM_104_IS_INOUT(C_BRAM_104_IS_INOUT),
        .C_BRAM_105_IS_INOUT(C_BRAM_105_IS_INOUT),
        .C_BRAM_106_IS_INOUT(C_BRAM_106_IS_INOUT),
        .C_BRAM_107_IS_INOUT(C_BRAM_107_IS_INOUT),
        .C_BRAM_108_IS_INOUT(C_BRAM_108_IS_INOUT),
        .C_BRAM_109_IS_INOUT(C_BRAM_109_IS_INOUT),
        .C_BRAM_110_IS_INOUT(C_BRAM_110_IS_INOUT),
        .C_BRAM_111_IS_INOUT(C_BRAM_111_IS_INOUT),
        .C_BRAM_112_IS_INOUT(C_BRAM_112_IS_INOUT),
        .C_BRAM_113_IS_INOUT(C_BRAM_113_IS_INOUT),
        .C_BRAM_114_IS_INOUT(C_BRAM_114_IS_INOUT),
        .C_BRAM_115_IS_INOUT(C_BRAM_115_IS_INOUT),
        .C_BRAM_116_IS_INOUT(C_BRAM_116_IS_INOUT),
        .C_BRAM_117_IS_INOUT(C_BRAM_117_IS_INOUT),
        .C_BRAM_118_IS_INOUT(C_BRAM_118_IS_INOUT),
        .C_BRAM_119_IS_INOUT(C_BRAM_119_IS_INOUT),
        .C_BRAM_120_IS_INOUT(C_BRAM_120_IS_INOUT),
        .C_BRAM_121_IS_INOUT(C_BRAM_121_IS_INOUT),
        .C_BRAM_122_IS_INOUT(C_BRAM_122_IS_INOUT),
        .C_BRAM_123_IS_INOUT(C_BRAM_123_IS_INOUT),
        .C_BRAM_124_IS_INOUT(C_BRAM_124_IS_INOUT),
        .C_BRAM_125_IS_INOUT(C_BRAM_125_IS_INOUT),
        .C_BRAM_126_IS_INOUT(C_BRAM_126_IS_INOUT),
        .C_BRAM_127_IS_INOUT(C_BRAM_127_IS_INOUT),
        .C_INPUT_BRAM_0_MB_DEPTH(C_INPUT_BRAM_0_MB_DEPTH),
        .C_INPUT_BRAM_1_MB_DEPTH(C_INPUT_BRAM_1_MB_DEPTH),
        .C_INPUT_BRAM_2_MB_DEPTH(C_INPUT_BRAM_2_MB_DEPTH),
        .C_INPUT_BRAM_3_MB_DEPTH(C_INPUT_BRAM_3_MB_DEPTH),
        .C_INPUT_BRAM_4_MB_DEPTH(C_INPUT_BRAM_4_MB_DEPTH),
        .C_INPUT_BRAM_5_MB_DEPTH(C_INPUT_BRAM_5_MB_DEPTH),
        .C_INPUT_BRAM_6_MB_DEPTH(C_INPUT_BRAM_6_MB_DEPTH),
        .C_INPUT_BRAM_7_MB_DEPTH(C_INPUT_BRAM_7_MB_DEPTH),
        .C_INPUT_BRAM_8_MB_DEPTH(C_INPUT_BRAM_8_MB_DEPTH),
        .C_INPUT_BRAM_9_MB_DEPTH(C_INPUT_BRAM_9_MB_DEPTH),
        .C_INPUT_BRAM_10_MB_DEPTH(C_INPUT_BRAM_10_MB_DEPTH),
        .C_INPUT_BRAM_11_MB_DEPTH(C_INPUT_BRAM_11_MB_DEPTH),
        .C_INPUT_BRAM_12_MB_DEPTH(C_INPUT_BRAM_12_MB_DEPTH),
        .C_INPUT_BRAM_13_MB_DEPTH(C_INPUT_BRAM_13_MB_DEPTH),
        .C_INPUT_BRAM_14_MB_DEPTH(C_INPUT_BRAM_14_MB_DEPTH),
        .C_INPUT_BRAM_15_MB_DEPTH(C_INPUT_BRAM_15_MB_DEPTH),
        .C_INPUT_BRAM_16_MB_DEPTH(C_INPUT_BRAM_16_MB_DEPTH),
        .C_INPUT_BRAM_17_MB_DEPTH(C_INPUT_BRAM_17_MB_DEPTH),
        .C_INPUT_BRAM_18_MB_DEPTH(C_INPUT_BRAM_18_MB_DEPTH),
        .C_INPUT_BRAM_19_MB_DEPTH(C_INPUT_BRAM_19_MB_DEPTH),
        .C_INPUT_BRAM_20_MB_DEPTH(C_INPUT_BRAM_20_MB_DEPTH),
        .C_INPUT_BRAM_21_MB_DEPTH(C_INPUT_BRAM_21_MB_DEPTH),
        .C_INPUT_BRAM_22_MB_DEPTH(C_INPUT_BRAM_22_MB_DEPTH),
        .C_INPUT_BRAM_23_MB_DEPTH(C_INPUT_BRAM_23_MB_DEPTH),
        .C_INPUT_BRAM_24_MB_DEPTH(C_INPUT_BRAM_24_MB_DEPTH),
        .C_INPUT_BRAM_25_MB_DEPTH(C_INPUT_BRAM_25_MB_DEPTH),
        .C_INPUT_BRAM_26_MB_DEPTH(C_INPUT_BRAM_26_MB_DEPTH),
        .C_INPUT_BRAM_27_MB_DEPTH(C_INPUT_BRAM_27_MB_DEPTH),
        .C_INPUT_BRAM_28_MB_DEPTH(C_INPUT_BRAM_28_MB_DEPTH),
        .C_INPUT_BRAM_29_MB_DEPTH(C_INPUT_BRAM_29_MB_DEPTH),
        .C_INPUT_BRAM_30_MB_DEPTH(C_INPUT_BRAM_30_MB_DEPTH),
        .C_INPUT_BRAM_31_MB_DEPTH(C_INPUT_BRAM_31_MB_DEPTH),
        .C_INPUT_BRAM_32_MB_DEPTH(C_INPUT_BRAM_32_MB_DEPTH),
        .C_INPUT_BRAM_33_MB_DEPTH(C_INPUT_BRAM_33_MB_DEPTH),
        .C_INPUT_BRAM_34_MB_DEPTH(C_INPUT_BRAM_34_MB_DEPTH),
        .C_INPUT_BRAM_35_MB_DEPTH(C_INPUT_BRAM_35_MB_DEPTH),
        .C_INPUT_BRAM_36_MB_DEPTH(C_INPUT_BRAM_36_MB_DEPTH),
        .C_INPUT_BRAM_37_MB_DEPTH(C_INPUT_BRAM_37_MB_DEPTH),
        .C_INPUT_BRAM_38_MB_DEPTH(C_INPUT_BRAM_38_MB_DEPTH),
        .C_INPUT_BRAM_39_MB_DEPTH(C_INPUT_BRAM_39_MB_DEPTH),
        .C_INPUT_BRAM_40_MB_DEPTH(C_INPUT_BRAM_40_MB_DEPTH),
        .C_INPUT_BRAM_41_MB_DEPTH(C_INPUT_BRAM_41_MB_DEPTH),
        .C_INPUT_BRAM_42_MB_DEPTH(C_INPUT_BRAM_42_MB_DEPTH),
        .C_INPUT_BRAM_43_MB_DEPTH(C_INPUT_BRAM_43_MB_DEPTH),
        .C_INPUT_BRAM_44_MB_DEPTH(C_INPUT_BRAM_44_MB_DEPTH),
        .C_INPUT_BRAM_45_MB_DEPTH(C_INPUT_BRAM_45_MB_DEPTH),
        .C_INPUT_BRAM_46_MB_DEPTH(C_INPUT_BRAM_46_MB_DEPTH),
        .C_INPUT_BRAM_47_MB_DEPTH(C_INPUT_BRAM_47_MB_DEPTH),
        .C_INPUT_BRAM_48_MB_DEPTH(C_INPUT_BRAM_48_MB_DEPTH),
        .C_INPUT_BRAM_49_MB_DEPTH(C_INPUT_BRAM_49_MB_DEPTH),
        .C_INPUT_BRAM_50_MB_DEPTH(C_INPUT_BRAM_50_MB_DEPTH),
        .C_INPUT_BRAM_51_MB_DEPTH(C_INPUT_BRAM_51_MB_DEPTH),
        .C_INPUT_BRAM_52_MB_DEPTH(C_INPUT_BRAM_52_MB_DEPTH),
        .C_INPUT_BRAM_53_MB_DEPTH(C_INPUT_BRAM_53_MB_DEPTH),
        .C_INPUT_BRAM_54_MB_DEPTH(C_INPUT_BRAM_54_MB_DEPTH),
        .C_INPUT_BRAM_55_MB_DEPTH(C_INPUT_BRAM_55_MB_DEPTH),
        .C_INPUT_BRAM_56_MB_DEPTH(C_INPUT_BRAM_56_MB_DEPTH),
        .C_INPUT_BRAM_57_MB_DEPTH(C_INPUT_BRAM_57_MB_DEPTH),
        .C_INPUT_BRAM_58_MB_DEPTH(C_INPUT_BRAM_58_MB_DEPTH),
        .C_INPUT_BRAM_59_MB_DEPTH(C_INPUT_BRAM_59_MB_DEPTH),
        .C_INPUT_BRAM_60_MB_DEPTH(C_INPUT_BRAM_60_MB_DEPTH),
        .C_INPUT_BRAM_61_MB_DEPTH(C_INPUT_BRAM_61_MB_DEPTH),
        .C_INPUT_BRAM_62_MB_DEPTH(C_INPUT_BRAM_62_MB_DEPTH),
        .C_INPUT_BRAM_63_MB_DEPTH(C_INPUT_BRAM_63_MB_DEPTH),
        .C_INPUT_BRAM_64_MB_DEPTH(C_INPUT_BRAM_64_MB_DEPTH),
        .C_INPUT_BRAM_65_MB_DEPTH(C_INPUT_BRAM_65_MB_DEPTH),
        .C_INPUT_BRAM_66_MB_DEPTH(C_INPUT_BRAM_66_MB_DEPTH),
        .C_INPUT_BRAM_67_MB_DEPTH(C_INPUT_BRAM_67_MB_DEPTH),
        .C_INPUT_BRAM_68_MB_DEPTH(C_INPUT_BRAM_68_MB_DEPTH),
        .C_INPUT_BRAM_69_MB_DEPTH(C_INPUT_BRAM_69_MB_DEPTH),
        .C_INPUT_BRAM_70_MB_DEPTH(C_INPUT_BRAM_70_MB_DEPTH),
        .C_INPUT_BRAM_71_MB_DEPTH(C_INPUT_BRAM_71_MB_DEPTH),
        .C_INPUT_BRAM_72_MB_DEPTH(C_INPUT_BRAM_72_MB_DEPTH),
        .C_INPUT_BRAM_73_MB_DEPTH(C_INPUT_BRAM_73_MB_DEPTH),
        .C_INPUT_BRAM_74_MB_DEPTH(C_INPUT_BRAM_74_MB_DEPTH),
        .C_INPUT_BRAM_75_MB_DEPTH(C_INPUT_BRAM_75_MB_DEPTH),
        .C_INPUT_BRAM_76_MB_DEPTH(C_INPUT_BRAM_76_MB_DEPTH),
        .C_INPUT_BRAM_77_MB_DEPTH(C_INPUT_BRAM_77_MB_DEPTH),
        .C_INPUT_BRAM_78_MB_DEPTH(C_INPUT_BRAM_78_MB_DEPTH),
        .C_INPUT_BRAM_79_MB_DEPTH(C_INPUT_BRAM_79_MB_DEPTH),
        .C_INPUT_BRAM_80_MB_DEPTH(C_INPUT_BRAM_80_MB_DEPTH),
        .C_INPUT_BRAM_81_MB_DEPTH(C_INPUT_BRAM_81_MB_DEPTH),
        .C_INPUT_BRAM_82_MB_DEPTH(C_INPUT_BRAM_82_MB_DEPTH),
        .C_INPUT_BRAM_83_MB_DEPTH(C_INPUT_BRAM_83_MB_DEPTH),
        .C_INPUT_BRAM_84_MB_DEPTH(C_INPUT_BRAM_84_MB_DEPTH),
        .C_INPUT_BRAM_85_MB_DEPTH(C_INPUT_BRAM_85_MB_DEPTH),
        .C_INPUT_BRAM_86_MB_DEPTH(C_INPUT_BRAM_86_MB_DEPTH),
        .C_INPUT_BRAM_87_MB_DEPTH(C_INPUT_BRAM_87_MB_DEPTH),
        .C_INPUT_BRAM_88_MB_DEPTH(C_INPUT_BRAM_88_MB_DEPTH),
        .C_INPUT_BRAM_89_MB_DEPTH(C_INPUT_BRAM_89_MB_DEPTH),
        .C_INPUT_BRAM_90_MB_DEPTH(C_INPUT_BRAM_90_MB_DEPTH),
        .C_INPUT_BRAM_91_MB_DEPTH(C_INPUT_BRAM_91_MB_DEPTH),
        .C_INPUT_BRAM_92_MB_DEPTH(C_INPUT_BRAM_92_MB_DEPTH),
        .C_INPUT_BRAM_93_MB_DEPTH(C_INPUT_BRAM_93_MB_DEPTH),
        .C_INPUT_BRAM_94_MB_DEPTH(C_INPUT_BRAM_94_MB_DEPTH),
        .C_INPUT_BRAM_95_MB_DEPTH(C_INPUT_BRAM_95_MB_DEPTH),
        .C_INPUT_BRAM_96_MB_DEPTH(C_INPUT_BRAM_96_MB_DEPTH),
        .C_INPUT_BRAM_97_MB_DEPTH(C_INPUT_BRAM_97_MB_DEPTH),
        .C_INPUT_BRAM_98_MB_DEPTH(C_INPUT_BRAM_98_MB_DEPTH),
        .C_INPUT_BRAM_99_MB_DEPTH(C_INPUT_BRAM_99_MB_DEPTH),
        .C_INPUT_BRAM_100_MB_DEPTH(C_INPUT_BRAM_100_MB_DEPTH),
        .C_INPUT_BRAM_101_MB_DEPTH(C_INPUT_BRAM_101_MB_DEPTH),
        .C_INPUT_BRAM_102_MB_DEPTH(C_INPUT_BRAM_102_MB_DEPTH),
        .C_INPUT_BRAM_103_MB_DEPTH(C_INPUT_BRAM_103_MB_DEPTH),
        .C_INPUT_BRAM_104_MB_DEPTH(C_INPUT_BRAM_104_MB_DEPTH),
        .C_INPUT_BRAM_105_MB_DEPTH(C_INPUT_BRAM_105_MB_DEPTH),
        .C_INPUT_BRAM_106_MB_DEPTH(C_INPUT_BRAM_106_MB_DEPTH),
        .C_INPUT_BRAM_107_MB_DEPTH(C_INPUT_BRAM_107_MB_DEPTH),
        .C_INPUT_BRAM_108_MB_DEPTH(C_INPUT_BRAM_108_MB_DEPTH),
        .C_INPUT_BRAM_109_MB_DEPTH(C_INPUT_BRAM_109_MB_DEPTH),
        .C_INPUT_BRAM_110_MB_DEPTH(C_INPUT_BRAM_110_MB_DEPTH),
        .C_INPUT_BRAM_111_MB_DEPTH(C_INPUT_BRAM_111_MB_DEPTH),
        .C_INPUT_BRAM_112_MB_DEPTH(C_INPUT_BRAM_112_MB_DEPTH),
        .C_INPUT_BRAM_113_MB_DEPTH(C_INPUT_BRAM_113_MB_DEPTH),
        .C_INPUT_BRAM_114_MB_DEPTH(C_INPUT_BRAM_114_MB_DEPTH),
        .C_INPUT_BRAM_115_MB_DEPTH(C_INPUT_BRAM_115_MB_DEPTH),
        .C_INPUT_BRAM_116_MB_DEPTH(C_INPUT_BRAM_116_MB_DEPTH),
        .C_INPUT_BRAM_117_MB_DEPTH(C_INPUT_BRAM_117_MB_DEPTH),
        .C_INPUT_BRAM_118_MB_DEPTH(C_INPUT_BRAM_118_MB_DEPTH),
        .C_INPUT_BRAM_119_MB_DEPTH(C_INPUT_BRAM_119_MB_DEPTH),
        .C_INPUT_BRAM_120_MB_DEPTH(C_INPUT_BRAM_120_MB_DEPTH),
        .C_INPUT_BRAM_121_MB_DEPTH(C_INPUT_BRAM_121_MB_DEPTH),
        .C_INPUT_BRAM_122_MB_DEPTH(C_INPUT_BRAM_122_MB_DEPTH),
        .C_INPUT_BRAM_123_MB_DEPTH(C_INPUT_BRAM_123_MB_DEPTH),
        .C_INPUT_BRAM_124_MB_DEPTH(C_INPUT_BRAM_124_MB_DEPTH),
        .C_INPUT_BRAM_125_MB_DEPTH(C_INPUT_BRAM_125_MB_DEPTH),
        .C_INPUT_BRAM_126_MB_DEPTH(C_INPUT_BRAM_126_MB_DEPTH),
        .C_INPUT_BRAM_127_MB_DEPTH(C_INPUT_BRAM_127_MB_DEPTH),
        .C_INPUT_BRAM_0_ADDR_WIDTH(C_INPUT_BRAM_0_ADDR_WIDTH),
        .C_INPUT_BRAM_1_ADDR_WIDTH(C_INPUT_BRAM_1_ADDR_WIDTH),
        .C_INPUT_BRAM_2_ADDR_WIDTH(C_INPUT_BRAM_2_ADDR_WIDTH),
        .C_INPUT_BRAM_3_ADDR_WIDTH(C_INPUT_BRAM_3_ADDR_WIDTH),
        .C_INPUT_BRAM_4_ADDR_WIDTH(C_INPUT_BRAM_4_ADDR_WIDTH),
        .C_INPUT_BRAM_5_ADDR_WIDTH(C_INPUT_BRAM_5_ADDR_WIDTH),
        .C_INPUT_BRAM_6_ADDR_WIDTH(C_INPUT_BRAM_6_ADDR_WIDTH),
        .C_INPUT_BRAM_7_ADDR_WIDTH(C_INPUT_BRAM_7_ADDR_WIDTH),
        .C_INPUT_BRAM_8_ADDR_WIDTH(C_INPUT_BRAM_8_ADDR_WIDTH),
        .C_INPUT_BRAM_9_ADDR_WIDTH(C_INPUT_BRAM_9_ADDR_WIDTH),
        .C_INPUT_BRAM_10_ADDR_WIDTH(C_INPUT_BRAM_10_ADDR_WIDTH),
        .C_INPUT_BRAM_11_ADDR_WIDTH(C_INPUT_BRAM_11_ADDR_WIDTH),
        .C_INPUT_BRAM_12_ADDR_WIDTH(C_INPUT_BRAM_12_ADDR_WIDTH),
        .C_INPUT_BRAM_13_ADDR_WIDTH(C_INPUT_BRAM_13_ADDR_WIDTH),
        .C_INPUT_BRAM_14_ADDR_WIDTH(C_INPUT_BRAM_14_ADDR_WIDTH),
        .C_INPUT_BRAM_15_ADDR_WIDTH(C_INPUT_BRAM_15_ADDR_WIDTH),
        .C_INPUT_BRAM_16_ADDR_WIDTH(C_INPUT_BRAM_16_ADDR_WIDTH),
        .C_INPUT_BRAM_17_ADDR_WIDTH(C_INPUT_BRAM_17_ADDR_WIDTH),
        .C_INPUT_BRAM_18_ADDR_WIDTH(C_INPUT_BRAM_18_ADDR_WIDTH),
        .C_INPUT_BRAM_19_ADDR_WIDTH(C_INPUT_BRAM_19_ADDR_WIDTH),
        .C_INPUT_BRAM_20_ADDR_WIDTH(C_INPUT_BRAM_20_ADDR_WIDTH),
        .C_INPUT_BRAM_21_ADDR_WIDTH(C_INPUT_BRAM_21_ADDR_WIDTH),
        .C_INPUT_BRAM_22_ADDR_WIDTH(C_INPUT_BRAM_22_ADDR_WIDTH),
        .C_INPUT_BRAM_23_ADDR_WIDTH(C_INPUT_BRAM_23_ADDR_WIDTH),
        .C_INPUT_BRAM_24_ADDR_WIDTH(C_INPUT_BRAM_24_ADDR_WIDTH),
        .C_INPUT_BRAM_25_ADDR_WIDTH(C_INPUT_BRAM_25_ADDR_WIDTH),
        .C_INPUT_BRAM_26_ADDR_WIDTH(C_INPUT_BRAM_26_ADDR_WIDTH),
        .C_INPUT_BRAM_27_ADDR_WIDTH(C_INPUT_BRAM_27_ADDR_WIDTH),
        .C_INPUT_BRAM_28_ADDR_WIDTH(C_INPUT_BRAM_28_ADDR_WIDTH),
        .C_INPUT_BRAM_29_ADDR_WIDTH(C_INPUT_BRAM_29_ADDR_WIDTH),
        .C_INPUT_BRAM_30_ADDR_WIDTH(C_INPUT_BRAM_30_ADDR_WIDTH),
        .C_INPUT_BRAM_31_ADDR_WIDTH(C_INPUT_BRAM_31_ADDR_WIDTH),
        .C_INPUT_BRAM_32_ADDR_WIDTH(C_INPUT_BRAM_32_ADDR_WIDTH),
        .C_INPUT_BRAM_33_ADDR_WIDTH(C_INPUT_BRAM_33_ADDR_WIDTH),
        .C_INPUT_BRAM_34_ADDR_WIDTH(C_INPUT_BRAM_34_ADDR_WIDTH),
        .C_INPUT_BRAM_35_ADDR_WIDTH(C_INPUT_BRAM_35_ADDR_WIDTH),
        .C_INPUT_BRAM_36_ADDR_WIDTH(C_INPUT_BRAM_36_ADDR_WIDTH),
        .C_INPUT_BRAM_37_ADDR_WIDTH(C_INPUT_BRAM_37_ADDR_WIDTH),
        .C_INPUT_BRAM_38_ADDR_WIDTH(C_INPUT_BRAM_38_ADDR_WIDTH),
        .C_INPUT_BRAM_39_ADDR_WIDTH(C_INPUT_BRAM_39_ADDR_WIDTH),
        .C_INPUT_BRAM_40_ADDR_WIDTH(C_INPUT_BRAM_40_ADDR_WIDTH),
        .C_INPUT_BRAM_41_ADDR_WIDTH(C_INPUT_BRAM_41_ADDR_WIDTH),
        .C_INPUT_BRAM_42_ADDR_WIDTH(C_INPUT_BRAM_42_ADDR_WIDTH),
        .C_INPUT_BRAM_43_ADDR_WIDTH(C_INPUT_BRAM_43_ADDR_WIDTH),
        .C_INPUT_BRAM_44_ADDR_WIDTH(C_INPUT_BRAM_44_ADDR_WIDTH),
        .C_INPUT_BRAM_45_ADDR_WIDTH(C_INPUT_BRAM_45_ADDR_WIDTH),
        .C_INPUT_BRAM_46_ADDR_WIDTH(C_INPUT_BRAM_46_ADDR_WIDTH),
        .C_INPUT_BRAM_47_ADDR_WIDTH(C_INPUT_BRAM_47_ADDR_WIDTH),
        .C_INPUT_BRAM_48_ADDR_WIDTH(C_INPUT_BRAM_48_ADDR_WIDTH),
        .C_INPUT_BRAM_49_ADDR_WIDTH(C_INPUT_BRAM_49_ADDR_WIDTH),
        .C_INPUT_BRAM_50_ADDR_WIDTH(C_INPUT_BRAM_50_ADDR_WIDTH),
        .C_INPUT_BRAM_51_ADDR_WIDTH(C_INPUT_BRAM_51_ADDR_WIDTH),
        .C_INPUT_BRAM_52_ADDR_WIDTH(C_INPUT_BRAM_52_ADDR_WIDTH),
        .C_INPUT_BRAM_53_ADDR_WIDTH(C_INPUT_BRAM_53_ADDR_WIDTH),
        .C_INPUT_BRAM_54_ADDR_WIDTH(C_INPUT_BRAM_54_ADDR_WIDTH),
        .C_INPUT_BRAM_55_ADDR_WIDTH(C_INPUT_BRAM_55_ADDR_WIDTH),
        .C_INPUT_BRAM_56_ADDR_WIDTH(C_INPUT_BRAM_56_ADDR_WIDTH),
        .C_INPUT_BRAM_57_ADDR_WIDTH(C_INPUT_BRAM_57_ADDR_WIDTH),
        .C_INPUT_BRAM_58_ADDR_WIDTH(C_INPUT_BRAM_58_ADDR_WIDTH),
        .C_INPUT_BRAM_59_ADDR_WIDTH(C_INPUT_BRAM_59_ADDR_WIDTH),
        .C_INPUT_BRAM_60_ADDR_WIDTH(C_INPUT_BRAM_60_ADDR_WIDTH),
        .C_INPUT_BRAM_61_ADDR_WIDTH(C_INPUT_BRAM_61_ADDR_WIDTH),
        .C_INPUT_BRAM_62_ADDR_WIDTH(C_INPUT_BRAM_62_ADDR_WIDTH),
        .C_INPUT_BRAM_63_ADDR_WIDTH(C_INPUT_BRAM_63_ADDR_WIDTH),
        .C_INPUT_BRAM_64_ADDR_WIDTH(C_INPUT_BRAM_64_ADDR_WIDTH),
        .C_INPUT_BRAM_65_ADDR_WIDTH(C_INPUT_BRAM_65_ADDR_WIDTH),
        .C_INPUT_BRAM_66_ADDR_WIDTH(C_INPUT_BRAM_66_ADDR_WIDTH),
        .C_INPUT_BRAM_67_ADDR_WIDTH(C_INPUT_BRAM_67_ADDR_WIDTH),
        .C_INPUT_BRAM_68_ADDR_WIDTH(C_INPUT_BRAM_68_ADDR_WIDTH),
        .C_INPUT_BRAM_69_ADDR_WIDTH(C_INPUT_BRAM_69_ADDR_WIDTH),
        .C_INPUT_BRAM_70_ADDR_WIDTH(C_INPUT_BRAM_70_ADDR_WIDTH),
        .C_INPUT_BRAM_71_ADDR_WIDTH(C_INPUT_BRAM_71_ADDR_WIDTH),
        .C_INPUT_BRAM_72_ADDR_WIDTH(C_INPUT_BRAM_72_ADDR_WIDTH),
        .C_INPUT_BRAM_73_ADDR_WIDTH(C_INPUT_BRAM_73_ADDR_WIDTH),
        .C_INPUT_BRAM_74_ADDR_WIDTH(C_INPUT_BRAM_74_ADDR_WIDTH),
        .C_INPUT_BRAM_75_ADDR_WIDTH(C_INPUT_BRAM_75_ADDR_WIDTH),
        .C_INPUT_BRAM_76_ADDR_WIDTH(C_INPUT_BRAM_76_ADDR_WIDTH),
        .C_INPUT_BRAM_77_ADDR_WIDTH(C_INPUT_BRAM_77_ADDR_WIDTH),
        .C_INPUT_BRAM_78_ADDR_WIDTH(C_INPUT_BRAM_78_ADDR_WIDTH),
        .C_INPUT_BRAM_79_ADDR_WIDTH(C_INPUT_BRAM_79_ADDR_WIDTH),
        .C_INPUT_BRAM_80_ADDR_WIDTH(C_INPUT_BRAM_80_ADDR_WIDTH),
        .C_INPUT_BRAM_81_ADDR_WIDTH(C_INPUT_BRAM_81_ADDR_WIDTH),
        .C_INPUT_BRAM_82_ADDR_WIDTH(C_INPUT_BRAM_82_ADDR_WIDTH),
        .C_INPUT_BRAM_83_ADDR_WIDTH(C_INPUT_BRAM_83_ADDR_WIDTH),
        .C_INPUT_BRAM_84_ADDR_WIDTH(C_INPUT_BRAM_84_ADDR_WIDTH),
        .C_INPUT_BRAM_85_ADDR_WIDTH(C_INPUT_BRAM_85_ADDR_WIDTH),
        .C_INPUT_BRAM_86_ADDR_WIDTH(C_INPUT_BRAM_86_ADDR_WIDTH),
        .C_INPUT_BRAM_87_ADDR_WIDTH(C_INPUT_BRAM_87_ADDR_WIDTH),
        .C_INPUT_BRAM_88_ADDR_WIDTH(C_INPUT_BRAM_88_ADDR_WIDTH),
        .C_INPUT_BRAM_89_ADDR_WIDTH(C_INPUT_BRAM_89_ADDR_WIDTH),
        .C_INPUT_BRAM_90_ADDR_WIDTH(C_INPUT_BRAM_90_ADDR_WIDTH),
        .C_INPUT_BRAM_91_ADDR_WIDTH(C_INPUT_BRAM_91_ADDR_WIDTH),
        .C_INPUT_BRAM_92_ADDR_WIDTH(C_INPUT_BRAM_92_ADDR_WIDTH),
        .C_INPUT_BRAM_93_ADDR_WIDTH(C_INPUT_BRAM_93_ADDR_WIDTH),
        .C_INPUT_BRAM_94_ADDR_WIDTH(C_INPUT_BRAM_94_ADDR_WIDTH),
        .C_INPUT_BRAM_95_ADDR_WIDTH(C_INPUT_BRAM_95_ADDR_WIDTH),
        .C_INPUT_BRAM_96_ADDR_WIDTH(C_INPUT_BRAM_96_ADDR_WIDTH),
        .C_INPUT_BRAM_97_ADDR_WIDTH(C_INPUT_BRAM_97_ADDR_WIDTH),
        .C_INPUT_BRAM_98_ADDR_WIDTH(C_INPUT_BRAM_98_ADDR_WIDTH),
        .C_INPUT_BRAM_99_ADDR_WIDTH(C_INPUT_BRAM_99_ADDR_WIDTH),
        .C_INPUT_BRAM_100_ADDR_WIDTH(C_INPUT_BRAM_100_ADDR_WIDTH),
        .C_INPUT_BRAM_101_ADDR_WIDTH(C_INPUT_BRAM_101_ADDR_WIDTH),
        .C_INPUT_BRAM_102_ADDR_WIDTH(C_INPUT_BRAM_102_ADDR_WIDTH),
        .C_INPUT_BRAM_103_ADDR_WIDTH(C_INPUT_BRAM_103_ADDR_WIDTH),
        .C_INPUT_BRAM_104_ADDR_WIDTH(C_INPUT_BRAM_104_ADDR_WIDTH),
        .C_INPUT_BRAM_105_ADDR_WIDTH(C_INPUT_BRAM_105_ADDR_WIDTH),
        .C_INPUT_BRAM_106_ADDR_WIDTH(C_INPUT_BRAM_106_ADDR_WIDTH),
        .C_INPUT_BRAM_107_ADDR_WIDTH(C_INPUT_BRAM_107_ADDR_WIDTH),
        .C_INPUT_BRAM_108_ADDR_WIDTH(C_INPUT_BRAM_108_ADDR_WIDTH),
        .C_INPUT_BRAM_109_ADDR_WIDTH(C_INPUT_BRAM_109_ADDR_WIDTH),
        .C_INPUT_BRAM_110_ADDR_WIDTH(C_INPUT_BRAM_110_ADDR_WIDTH),
        .C_INPUT_BRAM_111_ADDR_WIDTH(C_INPUT_BRAM_111_ADDR_WIDTH),
        .C_INPUT_BRAM_112_ADDR_WIDTH(C_INPUT_BRAM_112_ADDR_WIDTH),
        .C_INPUT_BRAM_113_ADDR_WIDTH(C_INPUT_BRAM_113_ADDR_WIDTH),
        .C_INPUT_BRAM_114_ADDR_WIDTH(C_INPUT_BRAM_114_ADDR_WIDTH),
        .C_INPUT_BRAM_115_ADDR_WIDTH(C_INPUT_BRAM_115_ADDR_WIDTH),
        .C_INPUT_BRAM_116_ADDR_WIDTH(C_INPUT_BRAM_116_ADDR_WIDTH),
        .C_INPUT_BRAM_117_ADDR_WIDTH(C_INPUT_BRAM_117_ADDR_WIDTH),
        .C_INPUT_BRAM_118_ADDR_WIDTH(C_INPUT_BRAM_118_ADDR_WIDTH),
        .C_INPUT_BRAM_119_ADDR_WIDTH(C_INPUT_BRAM_119_ADDR_WIDTH),
        .C_INPUT_BRAM_120_ADDR_WIDTH(C_INPUT_BRAM_120_ADDR_WIDTH),
        .C_INPUT_BRAM_121_ADDR_WIDTH(C_INPUT_BRAM_121_ADDR_WIDTH),
        .C_INPUT_BRAM_122_ADDR_WIDTH(C_INPUT_BRAM_122_ADDR_WIDTH),
        .C_INPUT_BRAM_123_ADDR_WIDTH(C_INPUT_BRAM_123_ADDR_WIDTH),
        .C_INPUT_BRAM_124_ADDR_WIDTH(C_INPUT_BRAM_124_ADDR_WIDTH),
        .C_INPUT_BRAM_125_ADDR_WIDTH(C_INPUT_BRAM_125_ADDR_WIDTH),
        .C_INPUT_BRAM_126_ADDR_WIDTH(C_INPUT_BRAM_126_ADDR_WIDTH),
        .C_INPUT_BRAM_127_ADDR_WIDTH(C_INPUT_BRAM_127_ADDR_WIDTH)
    ) in_bram_args_i (
        .acc_clk(aclk),
        .dm_clk(s_axi_aclk),
        .aresetn(s_axi_aresetn),
        .acc_rstn(resetn),
        .in_bram_allow_in(inbram_ctrl_allow),
        .in_bram_allow_out(outbram_ctrl_allow),
        .acc_start(ap_start_single),
        .acc_done(ap_done),
        .in_bram_ready(inbram_ctrl_ready),
        .inout_bram_ready(inoutbram_ctrl_ready),
        .s_axis_bram_0_tlast(s_axis_bram_0_tlast),
        .s_axis_bram_0_tvalid(s_axis_bram_0_tvalid),
        .s_axis_bram_0_tkeep(s_axis_bram_0_tkeep),
        .s_axis_bram_0_tstrb(s_axis_bram_0_tstrb),
        .s_axis_bram_0_tdata(s_axis_bram_0_tdata),
        .s_axis_bram_0_tready(s_axis_bram_0_tready),
        .ap_bram_0_addr0(ap_bram_iarg_0_addr0),
        .ap_bram_0_din0(ap_bram_iarg_0_din0),
        .ap_bram_0_dout0(ap_bram_iarg_0_dout0),
        .ap_bram_0_we0(ap_bram_iarg_0_we0),
        .ap_bram_0_en0(ap_bram_iarg_0_en0),
        .ap_bram_0_addr1(ap_bram_iarg_0_addr1),
        .ap_bram_0_din1(ap_bram_iarg_0_din1),
        .ap_bram_0_dout1(ap_bram_iarg_0_dout1),
        .ap_bram_0_we1(ap_bram_iarg_0_we1),
        .ap_bram_0_en1(ap_bram_iarg_0_en1),
        .s_axis_bram_1_tlast(s_axis_bram_1_tlast),
        .s_axis_bram_1_tvalid(s_axis_bram_1_tvalid),
        .s_axis_bram_1_tkeep(s_axis_bram_1_tkeep),
        .s_axis_bram_1_tstrb(s_axis_bram_1_tstrb),
        .s_axis_bram_1_tdata(s_axis_bram_1_tdata),
        .s_axis_bram_1_tready(s_axis_bram_1_tready),
        .ap_bram_1_addr0(ap_bram_iarg_1_addr0),
        .ap_bram_1_din0(ap_bram_iarg_1_din0),
        .ap_bram_1_dout0(ap_bram_iarg_1_dout0),
        .ap_bram_1_we0(ap_bram_iarg_1_we0),
        .ap_bram_1_en0(ap_bram_iarg_1_en0),
        .ap_bram_1_addr1(ap_bram_iarg_1_addr1),
        .ap_bram_1_din1(ap_bram_iarg_1_din1),
        .ap_bram_1_dout1(ap_bram_iarg_1_dout1),
        .ap_bram_1_we1(ap_bram_iarg_1_we1),
        .ap_bram_1_en1(ap_bram_iarg_1_en1),
        .s_axis_bram_2_tlast(s_axis_bram_2_tlast),
        .s_axis_bram_2_tvalid(s_axis_bram_2_tvalid),
        .s_axis_bram_2_tkeep(s_axis_bram_2_tkeep),
        .s_axis_bram_2_tstrb(s_axis_bram_2_tstrb),
        .s_axis_bram_2_tdata(s_axis_bram_2_tdata),
        .s_axis_bram_2_tready(s_axis_bram_2_tready),
        .ap_bram_2_addr0(ap_bram_iarg_2_addr0),
        .ap_bram_2_din0(ap_bram_iarg_2_din0),
        .ap_bram_2_dout0(ap_bram_iarg_2_dout0),
        .ap_bram_2_we0(ap_bram_iarg_2_we0),
        .ap_bram_2_en0(ap_bram_iarg_2_en0),
        .ap_bram_2_addr1(ap_bram_iarg_2_addr1),
        .ap_bram_2_din1(ap_bram_iarg_2_din1),
        .ap_bram_2_dout1(ap_bram_iarg_2_dout1),
        .ap_bram_2_we1(ap_bram_iarg_2_we1),
        .ap_bram_2_en1(ap_bram_iarg_2_en1),
        .s_axis_bram_3_tlast(s_axis_bram_3_tlast),
        .s_axis_bram_3_tvalid(s_axis_bram_3_tvalid),
        .s_axis_bram_3_tkeep(s_axis_bram_3_tkeep),
        .s_axis_bram_3_tstrb(s_axis_bram_3_tstrb),
        .s_axis_bram_3_tdata(s_axis_bram_3_tdata),
        .s_axis_bram_3_tready(s_axis_bram_3_tready),
        .ap_bram_3_addr0(ap_bram_iarg_3_addr0),
        .ap_bram_3_din0(ap_bram_iarg_3_din0),
        .ap_bram_3_dout0(ap_bram_iarg_3_dout0),
        .ap_bram_3_we0(ap_bram_iarg_3_we0),
        .ap_bram_3_en0(ap_bram_iarg_3_en0),
        .ap_bram_3_addr1(ap_bram_iarg_3_addr1),
        .ap_bram_3_din1(ap_bram_iarg_3_din1),
        .ap_bram_3_dout1(ap_bram_iarg_3_dout1),
        .ap_bram_3_we1(ap_bram_iarg_3_we1),
        .ap_bram_3_en1(ap_bram_iarg_3_en1),
        .s_axis_bram_4_tlast(s_axis_bram_4_tlast),
        .s_axis_bram_4_tvalid(s_axis_bram_4_tvalid),
        .s_axis_bram_4_tkeep(s_axis_bram_4_tkeep),
        .s_axis_bram_4_tstrb(s_axis_bram_4_tstrb),
        .s_axis_bram_4_tdata(s_axis_bram_4_tdata),
        .s_axis_bram_4_tready(s_axis_bram_4_tready),
        .ap_bram_4_addr0(ap_bram_iarg_4_addr0),
        .ap_bram_4_din0(ap_bram_iarg_4_din0),
        .ap_bram_4_dout0(ap_bram_iarg_4_dout0),
        .ap_bram_4_we0(ap_bram_iarg_4_we0),
        .ap_bram_4_en0(ap_bram_iarg_4_en0),
        .ap_bram_4_addr1(ap_bram_iarg_4_addr1),
        .ap_bram_4_din1(ap_bram_iarg_4_din1),
        .ap_bram_4_dout1(ap_bram_iarg_4_dout1),
        .ap_bram_4_we1(ap_bram_iarg_4_we1),
        .ap_bram_4_en1(ap_bram_iarg_4_en1),
        .s_axis_bram_5_tlast(s_axis_bram_5_tlast),
        .s_axis_bram_5_tvalid(s_axis_bram_5_tvalid),
        .s_axis_bram_5_tkeep(s_axis_bram_5_tkeep),
        .s_axis_bram_5_tstrb(s_axis_bram_5_tstrb),
        .s_axis_bram_5_tdata(s_axis_bram_5_tdata),
        .s_axis_bram_5_tready(s_axis_bram_5_tready),
        .ap_bram_5_addr0(ap_bram_iarg_5_addr0),
        .ap_bram_5_din0(ap_bram_iarg_5_din0),
        .ap_bram_5_dout0(ap_bram_iarg_5_dout0),
        .ap_bram_5_we0(ap_bram_iarg_5_we0),
        .ap_bram_5_en0(ap_bram_iarg_5_en0),
        .ap_bram_5_addr1(ap_bram_iarg_5_addr1),
        .ap_bram_5_din1(ap_bram_iarg_5_din1),
        .ap_bram_5_dout1(ap_bram_iarg_5_dout1),
        .ap_bram_5_we1(ap_bram_iarg_5_we1),
        .ap_bram_5_en1(ap_bram_iarg_5_en1),
        .s_axis_bram_6_tlast(s_axis_bram_6_tlast),
        .s_axis_bram_6_tvalid(s_axis_bram_6_tvalid),
        .s_axis_bram_6_tkeep(s_axis_bram_6_tkeep),
        .s_axis_bram_6_tstrb(s_axis_bram_6_tstrb),
        .s_axis_bram_6_tdata(s_axis_bram_6_tdata),
        .s_axis_bram_6_tready(s_axis_bram_6_tready),
        .ap_bram_6_addr0(ap_bram_iarg_6_addr0),
        .ap_bram_6_din0(ap_bram_iarg_6_din0),
        .ap_bram_6_dout0(ap_bram_iarg_6_dout0),
        .ap_bram_6_we0(ap_bram_iarg_6_we0),
        .ap_bram_6_en0(ap_bram_iarg_6_en0),
        .ap_bram_6_addr1(ap_bram_iarg_6_addr1),
        .ap_bram_6_din1(ap_bram_iarg_6_din1),
        .ap_bram_6_dout1(ap_bram_iarg_6_dout1),
        .ap_bram_6_we1(ap_bram_iarg_6_we1),
        .ap_bram_6_en1(ap_bram_iarg_6_en1),
        .s_axis_bram_7_tlast(s_axis_bram_7_tlast),
        .s_axis_bram_7_tvalid(s_axis_bram_7_tvalid),
        .s_axis_bram_7_tkeep(s_axis_bram_7_tkeep),
        .s_axis_bram_7_tstrb(s_axis_bram_7_tstrb),
        .s_axis_bram_7_tdata(s_axis_bram_7_tdata),
        .s_axis_bram_7_tready(s_axis_bram_7_tready),
        .ap_bram_7_addr0(ap_bram_iarg_7_addr0),
        .ap_bram_7_din0(ap_bram_iarg_7_din0),
        .ap_bram_7_dout0(ap_bram_iarg_7_dout0),
        .ap_bram_7_we0(ap_bram_iarg_7_we0),
        .ap_bram_7_en0(ap_bram_iarg_7_en0),
        .ap_bram_7_addr1(ap_bram_iarg_7_addr1),
        .ap_bram_7_din1(ap_bram_iarg_7_din1),
        .ap_bram_7_dout1(ap_bram_iarg_7_dout1),
        .ap_bram_7_we1(ap_bram_iarg_7_we1),
        .ap_bram_7_en1(ap_bram_iarg_7_en1),
        .s_axis_bram_8_tlast(s_axis_bram_8_tlast),
        .s_axis_bram_8_tvalid(s_axis_bram_8_tvalid),
        .s_axis_bram_8_tkeep(s_axis_bram_8_tkeep),
        .s_axis_bram_8_tstrb(s_axis_bram_8_tstrb),
        .s_axis_bram_8_tdata(s_axis_bram_8_tdata),
        .s_axis_bram_8_tready(s_axis_bram_8_tready),
        .ap_bram_8_addr0(ap_bram_iarg_8_addr0),
        .ap_bram_8_din0(ap_bram_iarg_8_din0),
        .ap_bram_8_dout0(ap_bram_iarg_8_dout0),
        .ap_bram_8_we0(ap_bram_iarg_8_we0),
        .ap_bram_8_en0(ap_bram_iarg_8_en0),
        .ap_bram_8_addr1(ap_bram_iarg_8_addr1),
        .ap_bram_8_din1(ap_bram_iarg_8_din1),
        .ap_bram_8_dout1(ap_bram_iarg_8_dout1),
        .ap_bram_8_we1(ap_bram_iarg_8_we1),
        .ap_bram_8_en1(ap_bram_iarg_8_en1),
        .s_axis_bram_9_tlast(s_axis_bram_9_tlast),
        .s_axis_bram_9_tvalid(s_axis_bram_9_tvalid),
        .s_axis_bram_9_tkeep(s_axis_bram_9_tkeep),
        .s_axis_bram_9_tstrb(s_axis_bram_9_tstrb),
        .s_axis_bram_9_tdata(s_axis_bram_9_tdata),
        .s_axis_bram_9_tready(s_axis_bram_9_tready),
        .ap_bram_9_addr0(ap_bram_iarg_9_addr0),
        .ap_bram_9_din0(ap_bram_iarg_9_din0),
        .ap_bram_9_dout0(ap_bram_iarg_9_dout0),
        .ap_bram_9_we0(ap_bram_iarg_9_we0),
        .ap_bram_9_en0(ap_bram_iarg_9_en0),
        .ap_bram_9_addr1(ap_bram_iarg_9_addr1),
        .ap_bram_9_din1(ap_bram_iarg_9_din1),
        .ap_bram_9_dout1(ap_bram_iarg_9_dout1),
        .ap_bram_9_we1(ap_bram_iarg_9_we1),
        .ap_bram_9_en1(ap_bram_iarg_9_en1),
        .s_axis_bram_10_tlast(s_axis_bram_10_tlast),
        .s_axis_bram_10_tvalid(s_axis_bram_10_tvalid),
        .s_axis_bram_10_tkeep(s_axis_bram_10_tkeep),
        .s_axis_bram_10_tstrb(s_axis_bram_10_tstrb),
        .s_axis_bram_10_tdata(s_axis_bram_10_tdata),
        .s_axis_bram_10_tready(s_axis_bram_10_tready),
        .ap_bram_10_addr0(ap_bram_iarg_10_addr0),
        .ap_bram_10_din0(ap_bram_iarg_10_din0),
        .ap_bram_10_dout0(ap_bram_iarg_10_dout0),
        .ap_bram_10_we0(ap_bram_iarg_10_we0),
        .ap_bram_10_en0(ap_bram_iarg_10_en0),
        .ap_bram_10_addr1(ap_bram_iarg_10_addr1),
        .ap_bram_10_din1(ap_bram_iarg_10_din1),
        .ap_bram_10_dout1(ap_bram_iarg_10_dout1),
        .ap_bram_10_we1(ap_bram_iarg_10_we1),
        .ap_bram_10_en1(ap_bram_iarg_10_en1),
        .s_axis_bram_11_tlast(s_axis_bram_11_tlast),
        .s_axis_bram_11_tvalid(s_axis_bram_11_tvalid),
        .s_axis_bram_11_tkeep(s_axis_bram_11_tkeep),
        .s_axis_bram_11_tstrb(s_axis_bram_11_tstrb),
        .s_axis_bram_11_tdata(s_axis_bram_11_tdata),
        .s_axis_bram_11_tready(s_axis_bram_11_tready),
        .ap_bram_11_addr0(ap_bram_iarg_11_addr0),
        .ap_bram_11_din0(ap_bram_iarg_11_din0),
        .ap_bram_11_dout0(ap_bram_iarg_11_dout0),
        .ap_bram_11_we0(ap_bram_iarg_11_we0),
        .ap_bram_11_en0(ap_bram_iarg_11_en0),
        .ap_bram_11_addr1(ap_bram_iarg_11_addr1),
        .ap_bram_11_din1(ap_bram_iarg_11_din1),
        .ap_bram_11_dout1(ap_bram_iarg_11_dout1),
        .ap_bram_11_we1(ap_bram_iarg_11_we1),
        .ap_bram_11_en1(ap_bram_iarg_11_en1),
        .s_axis_bram_12_tlast(s_axis_bram_12_tlast),
        .s_axis_bram_12_tvalid(s_axis_bram_12_tvalid),
        .s_axis_bram_12_tkeep(s_axis_bram_12_tkeep),
        .s_axis_bram_12_tstrb(s_axis_bram_12_tstrb),
        .s_axis_bram_12_tdata(s_axis_bram_12_tdata),
        .s_axis_bram_12_tready(s_axis_bram_12_tready),
        .ap_bram_12_addr0(ap_bram_iarg_12_addr0),
        .ap_bram_12_din0(ap_bram_iarg_12_din0),
        .ap_bram_12_dout0(ap_bram_iarg_12_dout0),
        .ap_bram_12_we0(ap_bram_iarg_12_we0),
        .ap_bram_12_en0(ap_bram_iarg_12_en0),
        .ap_bram_12_addr1(ap_bram_iarg_12_addr1),
        .ap_bram_12_din1(ap_bram_iarg_12_din1),
        .ap_bram_12_dout1(ap_bram_iarg_12_dout1),
        .ap_bram_12_we1(ap_bram_iarg_12_we1),
        .ap_bram_12_en1(ap_bram_iarg_12_en1),
        .s_axis_bram_13_tlast(s_axis_bram_13_tlast),
        .s_axis_bram_13_tvalid(s_axis_bram_13_tvalid),
        .s_axis_bram_13_tkeep(s_axis_bram_13_tkeep),
        .s_axis_bram_13_tstrb(s_axis_bram_13_tstrb),
        .s_axis_bram_13_tdata(s_axis_bram_13_tdata),
        .s_axis_bram_13_tready(s_axis_bram_13_tready),
        .ap_bram_13_addr0(ap_bram_iarg_13_addr0),
        .ap_bram_13_din0(ap_bram_iarg_13_din0),
        .ap_bram_13_dout0(ap_bram_iarg_13_dout0),
        .ap_bram_13_we0(ap_bram_iarg_13_we0),
        .ap_bram_13_en0(ap_bram_iarg_13_en0),
        .ap_bram_13_addr1(ap_bram_iarg_13_addr1),
        .ap_bram_13_din1(ap_bram_iarg_13_din1),
        .ap_bram_13_dout1(ap_bram_iarg_13_dout1),
        .ap_bram_13_we1(ap_bram_iarg_13_we1),
        .ap_bram_13_en1(ap_bram_iarg_13_en1),
        .s_axis_bram_14_tlast(s_axis_bram_14_tlast),
        .s_axis_bram_14_tvalid(s_axis_bram_14_tvalid),
        .s_axis_bram_14_tkeep(s_axis_bram_14_tkeep),
        .s_axis_bram_14_tstrb(s_axis_bram_14_tstrb),
        .s_axis_bram_14_tdata(s_axis_bram_14_tdata),
        .s_axis_bram_14_tready(s_axis_bram_14_tready),
        .ap_bram_14_addr0(ap_bram_iarg_14_addr0),
        .ap_bram_14_din0(ap_bram_iarg_14_din0),
        .ap_bram_14_dout0(ap_bram_iarg_14_dout0),
        .ap_bram_14_we0(ap_bram_iarg_14_we0),
        .ap_bram_14_en0(ap_bram_iarg_14_en0),
        .ap_bram_14_addr1(ap_bram_iarg_14_addr1),
        .ap_bram_14_din1(ap_bram_iarg_14_din1),
        .ap_bram_14_dout1(ap_bram_iarg_14_dout1),
        .ap_bram_14_we1(ap_bram_iarg_14_we1),
        .ap_bram_14_en1(ap_bram_iarg_14_en1),
        .s_axis_bram_15_tlast(s_axis_bram_15_tlast),
        .s_axis_bram_15_tvalid(s_axis_bram_15_tvalid),
        .s_axis_bram_15_tkeep(s_axis_bram_15_tkeep),
        .s_axis_bram_15_tstrb(s_axis_bram_15_tstrb),
        .s_axis_bram_15_tdata(s_axis_bram_15_tdata),
        .s_axis_bram_15_tready(s_axis_bram_15_tready),
        .ap_bram_15_addr0(ap_bram_iarg_15_addr0),
        .ap_bram_15_din0(ap_bram_iarg_15_din0),
        .ap_bram_15_dout0(ap_bram_iarg_15_dout0),
        .ap_bram_15_we0(ap_bram_iarg_15_we0),
        .ap_bram_15_en0(ap_bram_iarg_15_en0),
        .ap_bram_15_addr1(ap_bram_iarg_15_addr1),
        .ap_bram_15_din1(ap_bram_iarg_15_din1),
        .ap_bram_15_dout1(ap_bram_iarg_15_dout1),
        .ap_bram_15_we1(ap_bram_iarg_15_we1),
        .ap_bram_15_en1(ap_bram_iarg_15_en1),
        .s_axis_bram_16_tlast(s_axis_bram_16_tlast),
        .s_axis_bram_16_tvalid(s_axis_bram_16_tvalid),
        .s_axis_bram_16_tkeep(s_axis_bram_16_tkeep),
        .s_axis_bram_16_tstrb(s_axis_bram_16_tstrb),
        .s_axis_bram_16_tdata(s_axis_bram_16_tdata),
        .s_axis_bram_16_tready(s_axis_bram_16_tready),
        .ap_bram_16_addr0(ap_bram_iarg_16_addr0),
        .ap_bram_16_din0(ap_bram_iarg_16_din0),
        .ap_bram_16_dout0(ap_bram_iarg_16_dout0),
        .ap_bram_16_we0(ap_bram_iarg_16_we0),
        .ap_bram_16_en0(ap_bram_iarg_16_en0),
        .ap_bram_16_addr1(ap_bram_iarg_16_addr1),
        .ap_bram_16_din1(ap_bram_iarg_16_din1),
        .ap_bram_16_dout1(ap_bram_iarg_16_dout1),
        .ap_bram_16_we1(ap_bram_iarg_16_we1),
        .ap_bram_16_en1(ap_bram_iarg_16_en1),
        .s_axis_bram_17_tlast(s_axis_bram_17_tlast),
        .s_axis_bram_17_tvalid(s_axis_bram_17_tvalid),
        .s_axis_bram_17_tkeep(s_axis_bram_17_tkeep),
        .s_axis_bram_17_tstrb(s_axis_bram_17_tstrb),
        .s_axis_bram_17_tdata(s_axis_bram_17_tdata),
        .s_axis_bram_17_tready(s_axis_bram_17_tready),
        .ap_bram_17_addr0(ap_bram_iarg_17_addr0),
        .ap_bram_17_din0(ap_bram_iarg_17_din0),
        .ap_bram_17_dout0(ap_bram_iarg_17_dout0),
        .ap_bram_17_we0(ap_bram_iarg_17_we0),
        .ap_bram_17_en0(ap_bram_iarg_17_en0),
        .ap_bram_17_addr1(ap_bram_iarg_17_addr1),
        .ap_bram_17_din1(ap_bram_iarg_17_din1),
        .ap_bram_17_dout1(ap_bram_iarg_17_dout1),
        .ap_bram_17_we1(ap_bram_iarg_17_we1),
        .ap_bram_17_en1(ap_bram_iarg_17_en1),
        .s_axis_bram_18_tlast(s_axis_bram_18_tlast),
        .s_axis_bram_18_tvalid(s_axis_bram_18_tvalid),
        .s_axis_bram_18_tkeep(s_axis_bram_18_tkeep),
        .s_axis_bram_18_tstrb(s_axis_bram_18_tstrb),
        .s_axis_bram_18_tdata(s_axis_bram_18_tdata),
        .s_axis_bram_18_tready(s_axis_bram_18_tready),
        .ap_bram_18_addr0(ap_bram_iarg_18_addr0),
        .ap_bram_18_din0(ap_bram_iarg_18_din0),
        .ap_bram_18_dout0(ap_bram_iarg_18_dout0),
        .ap_bram_18_we0(ap_bram_iarg_18_we0),
        .ap_bram_18_en0(ap_bram_iarg_18_en0),
        .ap_bram_18_addr1(ap_bram_iarg_18_addr1),
        .ap_bram_18_din1(ap_bram_iarg_18_din1),
        .ap_bram_18_dout1(ap_bram_iarg_18_dout1),
        .ap_bram_18_we1(ap_bram_iarg_18_we1),
        .ap_bram_18_en1(ap_bram_iarg_18_en1),
        .s_axis_bram_19_tlast(s_axis_bram_19_tlast),
        .s_axis_bram_19_tvalid(s_axis_bram_19_tvalid),
        .s_axis_bram_19_tkeep(s_axis_bram_19_tkeep),
        .s_axis_bram_19_tstrb(s_axis_bram_19_tstrb),
        .s_axis_bram_19_tdata(s_axis_bram_19_tdata),
        .s_axis_bram_19_tready(s_axis_bram_19_tready),
        .ap_bram_19_addr0(ap_bram_iarg_19_addr0),
        .ap_bram_19_din0(ap_bram_iarg_19_din0),
        .ap_bram_19_dout0(ap_bram_iarg_19_dout0),
        .ap_bram_19_we0(ap_bram_iarg_19_we0),
        .ap_bram_19_en0(ap_bram_iarg_19_en0),
        .ap_bram_19_addr1(ap_bram_iarg_19_addr1),
        .ap_bram_19_din1(ap_bram_iarg_19_din1),
        .ap_bram_19_dout1(ap_bram_iarg_19_dout1),
        .ap_bram_19_we1(ap_bram_iarg_19_we1),
        .ap_bram_19_en1(ap_bram_iarg_19_en1),
        .s_axis_bram_20_tlast(s_axis_bram_20_tlast),
        .s_axis_bram_20_tvalid(s_axis_bram_20_tvalid),
        .s_axis_bram_20_tkeep(s_axis_bram_20_tkeep),
        .s_axis_bram_20_tstrb(s_axis_bram_20_tstrb),
        .s_axis_bram_20_tdata(s_axis_bram_20_tdata),
        .s_axis_bram_20_tready(s_axis_bram_20_tready),
        .ap_bram_20_addr0(ap_bram_iarg_20_addr0),
        .ap_bram_20_din0(ap_bram_iarg_20_din0),
        .ap_bram_20_dout0(ap_bram_iarg_20_dout0),
        .ap_bram_20_we0(ap_bram_iarg_20_we0),
        .ap_bram_20_en0(ap_bram_iarg_20_en0),
        .ap_bram_20_addr1(ap_bram_iarg_20_addr1),
        .ap_bram_20_din1(ap_bram_iarg_20_din1),
        .ap_bram_20_dout1(ap_bram_iarg_20_dout1),
        .ap_bram_20_we1(ap_bram_iarg_20_we1),
        .ap_bram_20_en1(ap_bram_iarg_20_en1),
        .s_axis_bram_21_tlast(s_axis_bram_21_tlast),
        .s_axis_bram_21_tvalid(s_axis_bram_21_tvalid),
        .s_axis_bram_21_tkeep(s_axis_bram_21_tkeep),
        .s_axis_bram_21_tstrb(s_axis_bram_21_tstrb),
        .s_axis_bram_21_tdata(s_axis_bram_21_tdata),
        .s_axis_bram_21_tready(s_axis_bram_21_tready),
        .ap_bram_21_addr0(ap_bram_iarg_21_addr0),
        .ap_bram_21_din0(ap_bram_iarg_21_din0),
        .ap_bram_21_dout0(ap_bram_iarg_21_dout0),
        .ap_bram_21_we0(ap_bram_iarg_21_we0),
        .ap_bram_21_en0(ap_bram_iarg_21_en0),
        .ap_bram_21_addr1(ap_bram_iarg_21_addr1),
        .ap_bram_21_din1(ap_bram_iarg_21_din1),
        .ap_bram_21_dout1(ap_bram_iarg_21_dout1),
        .ap_bram_21_we1(ap_bram_iarg_21_we1),
        .ap_bram_21_en1(ap_bram_iarg_21_en1),
        .s_axis_bram_22_tlast(s_axis_bram_22_tlast),
        .s_axis_bram_22_tvalid(s_axis_bram_22_tvalid),
        .s_axis_bram_22_tkeep(s_axis_bram_22_tkeep),
        .s_axis_bram_22_tstrb(s_axis_bram_22_tstrb),
        .s_axis_bram_22_tdata(s_axis_bram_22_tdata),
        .s_axis_bram_22_tready(s_axis_bram_22_tready),
        .ap_bram_22_addr0(ap_bram_iarg_22_addr0),
        .ap_bram_22_din0(ap_bram_iarg_22_din0),
        .ap_bram_22_dout0(ap_bram_iarg_22_dout0),
        .ap_bram_22_we0(ap_bram_iarg_22_we0),
        .ap_bram_22_en0(ap_bram_iarg_22_en0),
        .ap_bram_22_addr1(ap_bram_iarg_22_addr1),
        .ap_bram_22_din1(ap_bram_iarg_22_din1),
        .ap_bram_22_dout1(ap_bram_iarg_22_dout1),
        .ap_bram_22_we1(ap_bram_iarg_22_we1),
        .ap_bram_22_en1(ap_bram_iarg_22_en1),
        .s_axis_bram_23_tlast(s_axis_bram_23_tlast),
        .s_axis_bram_23_tvalid(s_axis_bram_23_tvalid),
        .s_axis_bram_23_tkeep(s_axis_bram_23_tkeep),
        .s_axis_bram_23_tstrb(s_axis_bram_23_tstrb),
        .s_axis_bram_23_tdata(s_axis_bram_23_tdata),
        .s_axis_bram_23_tready(s_axis_bram_23_tready),
        .ap_bram_23_addr0(ap_bram_iarg_23_addr0),
        .ap_bram_23_din0(ap_bram_iarg_23_din0),
        .ap_bram_23_dout0(ap_bram_iarg_23_dout0),
        .ap_bram_23_we0(ap_bram_iarg_23_we0),
        .ap_bram_23_en0(ap_bram_iarg_23_en0),
        .ap_bram_23_addr1(ap_bram_iarg_23_addr1),
        .ap_bram_23_din1(ap_bram_iarg_23_din1),
        .ap_bram_23_dout1(ap_bram_iarg_23_dout1),
        .ap_bram_23_we1(ap_bram_iarg_23_we1),
        .ap_bram_23_en1(ap_bram_iarg_23_en1),
        .s_axis_bram_24_tlast(s_axis_bram_24_tlast),
        .s_axis_bram_24_tvalid(s_axis_bram_24_tvalid),
        .s_axis_bram_24_tkeep(s_axis_bram_24_tkeep),
        .s_axis_bram_24_tstrb(s_axis_bram_24_tstrb),
        .s_axis_bram_24_tdata(s_axis_bram_24_tdata),
        .s_axis_bram_24_tready(s_axis_bram_24_tready),
        .ap_bram_24_addr0(ap_bram_iarg_24_addr0),
        .ap_bram_24_din0(ap_bram_iarg_24_din0),
        .ap_bram_24_dout0(ap_bram_iarg_24_dout0),
        .ap_bram_24_we0(ap_bram_iarg_24_we0),
        .ap_bram_24_en0(ap_bram_iarg_24_en0),
        .ap_bram_24_addr1(ap_bram_iarg_24_addr1),
        .ap_bram_24_din1(ap_bram_iarg_24_din1),
        .ap_bram_24_dout1(ap_bram_iarg_24_dout1),
        .ap_bram_24_we1(ap_bram_iarg_24_we1),
        .ap_bram_24_en1(ap_bram_iarg_24_en1),
        .s_axis_bram_25_tlast(s_axis_bram_25_tlast),
        .s_axis_bram_25_tvalid(s_axis_bram_25_tvalid),
        .s_axis_bram_25_tkeep(s_axis_bram_25_tkeep),
        .s_axis_bram_25_tstrb(s_axis_bram_25_tstrb),
        .s_axis_bram_25_tdata(s_axis_bram_25_tdata),
        .s_axis_bram_25_tready(s_axis_bram_25_tready),
        .ap_bram_25_addr0(ap_bram_iarg_25_addr0),
        .ap_bram_25_din0(ap_bram_iarg_25_din0),
        .ap_bram_25_dout0(ap_bram_iarg_25_dout0),
        .ap_bram_25_we0(ap_bram_iarg_25_we0),
        .ap_bram_25_en0(ap_bram_iarg_25_en0),
        .ap_bram_25_addr1(ap_bram_iarg_25_addr1),
        .ap_bram_25_din1(ap_bram_iarg_25_din1),
        .ap_bram_25_dout1(ap_bram_iarg_25_dout1),
        .ap_bram_25_we1(ap_bram_iarg_25_we1),
        .ap_bram_25_en1(ap_bram_iarg_25_en1),
        .s_axis_bram_26_tlast(s_axis_bram_26_tlast),
        .s_axis_bram_26_tvalid(s_axis_bram_26_tvalid),
        .s_axis_bram_26_tkeep(s_axis_bram_26_tkeep),
        .s_axis_bram_26_tstrb(s_axis_bram_26_tstrb),
        .s_axis_bram_26_tdata(s_axis_bram_26_tdata),
        .s_axis_bram_26_tready(s_axis_bram_26_tready),
        .ap_bram_26_addr0(ap_bram_iarg_26_addr0),
        .ap_bram_26_din0(ap_bram_iarg_26_din0),
        .ap_bram_26_dout0(ap_bram_iarg_26_dout0),
        .ap_bram_26_we0(ap_bram_iarg_26_we0),
        .ap_bram_26_en0(ap_bram_iarg_26_en0),
        .ap_bram_26_addr1(ap_bram_iarg_26_addr1),
        .ap_bram_26_din1(ap_bram_iarg_26_din1),
        .ap_bram_26_dout1(ap_bram_iarg_26_dout1),
        .ap_bram_26_we1(ap_bram_iarg_26_we1),
        .ap_bram_26_en1(ap_bram_iarg_26_en1),
        .s_axis_bram_27_tlast(s_axis_bram_27_tlast),
        .s_axis_bram_27_tvalid(s_axis_bram_27_tvalid),
        .s_axis_bram_27_tkeep(s_axis_bram_27_tkeep),
        .s_axis_bram_27_tstrb(s_axis_bram_27_tstrb),
        .s_axis_bram_27_tdata(s_axis_bram_27_tdata),
        .s_axis_bram_27_tready(s_axis_bram_27_tready),
        .ap_bram_27_addr0(ap_bram_iarg_27_addr0),
        .ap_bram_27_din0(ap_bram_iarg_27_din0),
        .ap_bram_27_dout0(ap_bram_iarg_27_dout0),
        .ap_bram_27_we0(ap_bram_iarg_27_we0),
        .ap_bram_27_en0(ap_bram_iarg_27_en0),
        .ap_bram_27_addr1(ap_bram_iarg_27_addr1),
        .ap_bram_27_din1(ap_bram_iarg_27_din1),
        .ap_bram_27_dout1(ap_bram_iarg_27_dout1),
        .ap_bram_27_we1(ap_bram_iarg_27_we1),
        .ap_bram_27_en1(ap_bram_iarg_27_en1),
        .s_axis_bram_28_tlast(s_axis_bram_28_tlast),
        .s_axis_bram_28_tvalid(s_axis_bram_28_tvalid),
        .s_axis_bram_28_tkeep(s_axis_bram_28_tkeep),
        .s_axis_bram_28_tstrb(s_axis_bram_28_tstrb),
        .s_axis_bram_28_tdata(s_axis_bram_28_tdata),
        .s_axis_bram_28_tready(s_axis_bram_28_tready),
        .ap_bram_28_addr0(ap_bram_iarg_28_addr0),
        .ap_bram_28_din0(ap_bram_iarg_28_din0),
        .ap_bram_28_dout0(ap_bram_iarg_28_dout0),
        .ap_bram_28_we0(ap_bram_iarg_28_we0),
        .ap_bram_28_en0(ap_bram_iarg_28_en0),
        .ap_bram_28_addr1(ap_bram_iarg_28_addr1),
        .ap_bram_28_din1(ap_bram_iarg_28_din1),
        .ap_bram_28_dout1(ap_bram_iarg_28_dout1),
        .ap_bram_28_we1(ap_bram_iarg_28_we1),
        .ap_bram_28_en1(ap_bram_iarg_28_en1),
        .s_axis_bram_29_tlast(s_axis_bram_29_tlast),
        .s_axis_bram_29_tvalid(s_axis_bram_29_tvalid),
        .s_axis_bram_29_tkeep(s_axis_bram_29_tkeep),
        .s_axis_bram_29_tstrb(s_axis_bram_29_tstrb),
        .s_axis_bram_29_tdata(s_axis_bram_29_tdata),
        .s_axis_bram_29_tready(s_axis_bram_29_tready),
        .ap_bram_29_addr0(ap_bram_iarg_29_addr0),
        .ap_bram_29_din0(ap_bram_iarg_29_din0),
        .ap_bram_29_dout0(ap_bram_iarg_29_dout0),
        .ap_bram_29_we0(ap_bram_iarg_29_we0),
        .ap_bram_29_en0(ap_bram_iarg_29_en0),
        .ap_bram_29_addr1(ap_bram_iarg_29_addr1),
        .ap_bram_29_din1(ap_bram_iarg_29_din1),
        .ap_bram_29_dout1(ap_bram_iarg_29_dout1),
        .ap_bram_29_we1(ap_bram_iarg_29_we1),
        .ap_bram_29_en1(ap_bram_iarg_29_en1),
        .s_axis_bram_30_tlast(s_axis_bram_30_tlast),
        .s_axis_bram_30_tvalid(s_axis_bram_30_tvalid),
        .s_axis_bram_30_tkeep(s_axis_bram_30_tkeep),
        .s_axis_bram_30_tstrb(s_axis_bram_30_tstrb),
        .s_axis_bram_30_tdata(s_axis_bram_30_tdata),
        .s_axis_bram_30_tready(s_axis_bram_30_tready),
        .ap_bram_30_addr0(ap_bram_iarg_30_addr0),
        .ap_bram_30_din0(ap_bram_iarg_30_din0),
        .ap_bram_30_dout0(ap_bram_iarg_30_dout0),
        .ap_bram_30_we0(ap_bram_iarg_30_we0),
        .ap_bram_30_en0(ap_bram_iarg_30_en0),
        .ap_bram_30_addr1(ap_bram_iarg_30_addr1),
        .ap_bram_30_din1(ap_bram_iarg_30_din1),
        .ap_bram_30_dout1(ap_bram_iarg_30_dout1),
        .ap_bram_30_we1(ap_bram_iarg_30_we1),
        .ap_bram_30_en1(ap_bram_iarg_30_en1),
        .s_axis_bram_31_tlast(s_axis_bram_31_tlast),
        .s_axis_bram_31_tvalid(s_axis_bram_31_tvalid),
        .s_axis_bram_31_tkeep(s_axis_bram_31_tkeep),
        .s_axis_bram_31_tstrb(s_axis_bram_31_tstrb),
        .s_axis_bram_31_tdata(s_axis_bram_31_tdata),
        .s_axis_bram_31_tready(s_axis_bram_31_tready),
        .ap_bram_31_addr0(ap_bram_iarg_31_addr0),
        .ap_bram_31_din0(ap_bram_iarg_31_din0),
        .ap_bram_31_dout0(ap_bram_iarg_31_dout0),
        .ap_bram_31_we0(ap_bram_iarg_31_we0),
        .ap_bram_31_en0(ap_bram_iarg_31_en0),
        .ap_bram_31_addr1(ap_bram_iarg_31_addr1),
        .ap_bram_31_din1(ap_bram_iarg_31_din1),
        .ap_bram_31_dout1(ap_bram_iarg_31_dout1),
        .ap_bram_31_we1(ap_bram_iarg_31_we1),
        .ap_bram_31_en1(ap_bram_iarg_31_en1),
        .s_axis_bram_32_tlast(s_axis_bram_32_tlast),
        .s_axis_bram_32_tvalid(s_axis_bram_32_tvalid),
        .s_axis_bram_32_tkeep(s_axis_bram_32_tkeep),
        .s_axis_bram_32_tstrb(s_axis_bram_32_tstrb),
        .s_axis_bram_32_tdata(s_axis_bram_32_tdata),
        .s_axis_bram_32_tready(s_axis_bram_32_tready),
        .ap_bram_32_addr0(ap_bram_iarg_32_addr0),
        .ap_bram_32_din0(ap_bram_iarg_32_din0),
        .ap_bram_32_dout0(ap_bram_iarg_32_dout0),
        .ap_bram_32_we0(ap_bram_iarg_32_we0),
        .ap_bram_32_en0(ap_bram_iarg_32_en0),
        .ap_bram_32_addr1(ap_bram_iarg_32_addr1),
        .ap_bram_32_din1(ap_bram_iarg_32_din1),
        .ap_bram_32_dout1(ap_bram_iarg_32_dout1),
        .ap_bram_32_we1(ap_bram_iarg_32_we1),
        .ap_bram_32_en1(ap_bram_iarg_32_en1),
        .s_axis_bram_33_tlast(s_axis_bram_33_tlast),
        .s_axis_bram_33_tvalid(s_axis_bram_33_tvalid),
        .s_axis_bram_33_tkeep(s_axis_bram_33_tkeep),
        .s_axis_bram_33_tstrb(s_axis_bram_33_tstrb),
        .s_axis_bram_33_tdata(s_axis_bram_33_tdata),
        .s_axis_bram_33_tready(s_axis_bram_33_tready),
        .ap_bram_33_addr0(ap_bram_iarg_33_addr0),
        .ap_bram_33_din0(ap_bram_iarg_33_din0),
        .ap_bram_33_dout0(ap_bram_iarg_33_dout0),
        .ap_bram_33_we0(ap_bram_iarg_33_we0),
        .ap_bram_33_en0(ap_bram_iarg_33_en0),
        .ap_bram_33_addr1(ap_bram_iarg_33_addr1),
        .ap_bram_33_din1(ap_bram_iarg_33_din1),
        .ap_bram_33_dout1(ap_bram_iarg_33_dout1),
        .ap_bram_33_we1(ap_bram_iarg_33_we1),
        .ap_bram_33_en1(ap_bram_iarg_33_en1),
        .s_axis_bram_34_tlast(s_axis_bram_34_tlast),
        .s_axis_bram_34_tvalid(s_axis_bram_34_tvalid),
        .s_axis_bram_34_tkeep(s_axis_bram_34_tkeep),
        .s_axis_bram_34_tstrb(s_axis_bram_34_tstrb),
        .s_axis_bram_34_tdata(s_axis_bram_34_tdata),
        .s_axis_bram_34_tready(s_axis_bram_34_tready),
        .ap_bram_34_addr0(ap_bram_iarg_34_addr0),
        .ap_bram_34_din0(ap_bram_iarg_34_din0),
        .ap_bram_34_dout0(ap_bram_iarg_34_dout0),
        .ap_bram_34_we0(ap_bram_iarg_34_we0),
        .ap_bram_34_en0(ap_bram_iarg_34_en0),
        .ap_bram_34_addr1(ap_bram_iarg_34_addr1),
        .ap_bram_34_din1(ap_bram_iarg_34_din1),
        .ap_bram_34_dout1(ap_bram_iarg_34_dout1),
        .ap_bram_34_we1(ap_bram_iarg_34_we1),
        .ap_bram_34_en1(ap_bram_iarg_34_en1),
        .s_axis_bram_35_tlast(s_axis_bram_35_tlast),
        .s_axis_bram_35_tvalid(s_axis_bram_35_tvalid),
        .s_axis_bram_35_tkeep(s_axis_bram_35_tkeep),
        .s_axis_bram_35_tstrb(s_axis_bram_35_tstrb),
        .s_axis_bram_35_tdata(s_axis_bram_35_tdata),
        .s_axis_bram_35_tready(s_axis_bram_35_tready),
        .ap_bram_35_addr0(ap_bram_iarg_35_addr0),
        .ap_bram_35_din0(ap_bram_iarg_35_din0),
        .ap_bram_35_dout0(ap_bram_iarg_35_dout0),
        .ap_bram_35_we0(ap_bram_iarg_35_we0),
        .ap_bram_35_en0(ap_bram_iarg_35_en0),
        .ap_bram_35_addr1(ap_bram_iarg_35_addr1),
        .ap_bram_35_din1(ap_bram_iarg_35_din1),
        .ap_bram_35_dout1(ap_bram_iarg_35_dout1),
        .ap_bram_35_we1(ap_bram_iarg_35_we1),
        .ap_bram_35_en1(ap_bram_iarg_35_en1),
        .s_axis_bram_36_tlast(s_axis_bram_36_tlast),
        .s_axis_bram_36_tvalid(s_axis_bram_36_tvalid),
        .s_axis_bram_36_tkeep(s_axis_bram_36_tkeep),
        .s_axis_bram_36_tstrb(s_axis_bram_36_tstrb),
        .s_axis_bram_36_tdata(s_axis_bram_36_tdata),
        .s_axis_bram_36_tready(s_axis_bram_36_tready),
        .ap_bram_36_addr0(ap_bram_iarg_36_addr0),
        .ap_bram_36_din0(ap_bram_iarg_36_din0),
        .ap_bram_36_dout0(ap_bram_iarg_36_dout0),
        .ap_bram_36_we0(ap_bram_iarg_36_we0),
        .ap_bram_36_en0(ap_bram_iarg_36_en0),
        .ap_bram_36_addr1(ap_bram_iarg_36_addr1),
        .ap_bram_36_din1(ap_bram_iarg_36_din1),
        .ap_bram_36_dout1(ap_bram_iarg_36_dout1),
        .ap_bram_36_we1(ap_bram_iarg_36_we1),
        .ap_bram_36_en1(ap_bram_iarg_36_en1),
        .s_axis_bram_37_tlast(s_axis_bram_37_tlast),
        .s_axis_bram_37_tvalid(s_axis_bram_37_tvalid),
        .s_axis_bram_37_tkeep(s_axis_bram_37_tkeep),
        .s_axis_bram_37_tstrb(s_axis_bram_37_tstrb),
        .s_axis_bram_37_tdata(s_axis_bram_37_tdata),
        .s_axis_bram_37_tready(s_axis_bram_37_tready),
        .ap_bram_37_addr0(ap_bram_iarg_37_addr0),
        .ap_bram_37_din0(ap_bram_iarg_37_din0),
        .ap_bram_37_dout0(ap_bram_iarg_37_dout0),
        .ap_bram_37_we0(ap_bram_iarg_37_we0),
        .ap_bram_37_en0(ap_bram_iarg_37_en0),
        .ap_bram_37_addr1(ap_bram_iarg_37_addr1),
        .ap_bram_37_din1(ap_bram_iarg_37_din1),
        .ap_bram_37_dout1(ap_bram_iarg_37_dout1),
        .ap_bram_37_we1(ap_bram_iarg_37_we1),
        .ap_bram_37_en1(ap_bram_iarg_37_en1),
        .s_axis_bram_38_tlast(s_axis_bram_38_tlast),
        .s_axis_bram_38_tvalid(s_axis_bram_38_tvalid),
        .s_axis_bram_38_tkeep(s_axis_bram_38_tkeep),
        .s_axis_bram_38_tstrb(s_axis_bram_38_tstrb),
        .s_axis_bram_38_tdata(s_axis_bram_38_tdata),
        .s_axis_bram_38_tready(s_axis_bram_38_tready),
        .ap_bram_38_addr0(ap_bram_iarg_38_addr0),
        .ap_bram_38_din0(ap_bram_iarg_38_din0),
        .ap_bram_38_dout0(ap_bram_iarg_38_dout0),
        .ap_bram_38_we0(ap_bram_iarg_38_we0),
        .ap_bram_38_en0(ap_bram_iarg_38_en0),
        .ap_bram_38_addr1(ap_bram_iarg_38_addr1),
        .ap_bram_38_din1(ap_bram_iarg_38_din1),
        .ap_bram_38_dout1(ap_bram_iarg_38_dout1),
        .ap_bram_38_we1(ap_bram_iarg_38_we1),
        .ap_bram_38_en1(ap_bram_iarg_38_en1),
        .s_axis_bram_39_tlast(s_axis_bram_39_tlast),
        .s_axis_bram_39_tvalid(s_axis_bram_39_tvalid),
        .s_axis_bram_39_tkeep(s_axis_bram_39_tkeep),
        .s_axis_bram_39_tstrb(s_axis_bram_39_tstrb),
        .s_axis_bram_39_tdata(s_axis_bram_39_tdata),
        .s_axis_bram_39_tready(s_axis_bram_39_tready),
        .ap_bram_39_addr0(ap_bram_iarg_39_addr0),
        .ap_bram_39_din0(ap_bram_iarg_39_din0),
        .ap_bram_39_dout0(ap_bram_iarg_39_dout0),
        .ap_bram_39_we0(ap_bram_iarg_39_we0),
        .ap_bram_39_en0(ap_bram_iarg_39_en0),
        .ap_bram_39_addr1(ap_bram_iarg_39_addr1),
        .ap_bram_39_din1(ap_bram_iarg_39_din1),
        .ap_bram_39_dout1(ap_bram_iarg_39_dout1),
        .ap_bram_39_we1(ap_bram_iarg_39_we1),
        .ap_bram_39_en1(ap_bram_iarg_39_en1),
        .s_axis_bram_40_tlast(s_axis_bram_40_tlast),
        .s_axis_bram_40_tvalid(s_axis_bram_40_tvalid),
        .s_axis_bram_40_tkeep(s_axis_bram_40_tkeep),
        .s_axis_bram_40_tstrb(s_axis_bram_40_tstrb),
        .s_axis_bram_40_tdata(s_axis_bram_40_tdata),
        .s_axis_bram_40_tready(s_axis_bram_40_tready),
        .ap_bram_40_addr0(ap_bram_iarg_40_addr0),
        .ap_bram_40_din0(ap_bram_iarg_40_din0),
        .ap_bram_40_dout0(ap_bram_iarg_40_dout0),
        .ap_bram_40_we0(ap_bram_iarg_40_we0),
        .ap_bram_40_en0(ap_bram_iarg_40_en0),
        .ap_bram_40_addr1(ap_bram_iarg_40_addr1),
        .ap_bram_40_din1(ap_bram_iarg_40_din1),
        .ap_bram_40_dout1(ap_bram_iarg_40_dout1),
        .ap_bram_40_we1(ap_bram_iarg_40_we1),
        .ap_bram_40_en1(ap_bram_iarg_40_en1),
        .s_axis_bram_41_tlast(s_axis_bram_41_tlast),
        .s_axis_bram_41_tvalid(s_axis_bram_41_tvalid),
        .s_axis_bram_41_tkeep(s_axis_bram_41_tkeep),
        .s_axis_bram_41_tstrb(s_axis_bram_41_tstrb),
        .s_axis_bram_41_tdata(s_axis_bram_41_tdata),
        .s_axis_bram_41_tready(s_axis_bram_41_tready),
        .ap_bram_41_addr0(ap_bram_iarg_41_addr0),
        .ap_bram_41_din0(ap_bram_iarg_41_din0),
        .ap_bram_41_dout0(ap_bram_iarg_41_dout0),
        .ap_bram_41_we0(ap_bram_iarg_41_we0),
        .ap_bram_41_en0(ap_bram_iarg_41_en0),
        .ap_bram_41_addr1(ap_bram_iarg_41_addr1),
        .ap_bram_41_din1(ap_bram_iarg_41_din1),
        .ap_bram_41_dout1(ap_bram_iarg_41_dout1),
        .ap_bram_41_we1(ap_bram_iarg_41_we1),
        .ap_bram_41_en1(ap_bram_iarg_41_en1),
        .s_axis_bram_42_tlast(s_axis_bram_42_tlast),
        .s_axis_bram_42_tvalid(s_axis_bram_42_tvalid),
        .s_axis_bram_42_tkeep(s_axis_bram_42_tkeep),
        .s_axis_bram_42_tstrb(s_axis_bram_42_tstrb),
        .s_axis_bram_42_tdata(s_axis_bram_42_tdata),
        .s_axis_bram_42_tready(s_axis_bram_42_tready),
        .ap_bram_42_addr0(ap_bram_iarg_42_addr0),
        .ap_bram_42_din0(ap_bram_iarg_42_din0),
        .ap_bram_42_dout0(ap_bram_iarg_42_dout0),
        .ap_bram_42_we0(ap_bram_iarg_42_we0),
        .ap_bram_42_en0(ap_bram_iarg_42_en0),
        .ap_bram_42_addr1(ap_bram_iarg_42_addr1),
        .ap_bram_42_din1(ap_bram_iarg_42_din1),
        .ap_bram_42_dout1(ap_bram_iarg_42_dout1),
        .ap_bram_42_we1(ap_bram_iarg_42_we1),
        .ap_bram_42_en1(ap_bram_iarg_42_en1),
        .s_axis_bram_43_tlast(s_axis_bram_43_tlast),
        .s_axis_bram_43_tvalid(s_axis_bram_43_tvalid),
        .s_axis_bram_43_tkeep(s_axis_bram_43_tkeep),
        .s_axis_bram_43_tstrb(s_axis_bram_43_tstrb),
        .s_axis_bram_43_tdata(s_axis_bram_43_tdata),
        .s_axis_bram_43_tready(s_axis_bram_43_tready),
        .ap_bram_43_addr0(ap_bram_iarg_43_addr0),
        .ap_bram_43_din0(ap_bram_iarg_43_din0),
        .ap_bram_43_dout0(ap_bram_iarg_43_dout0),
        .ap_bram_43_we0(ap_bram_iarg_43_we0),
        .ap_bram_43_en0(ap_bram_iarg_43_en0),
        .ap_bram_43_addr1(ap_bram_iarg_43_addr1),
        .ap_bram_43_din1(ap_bram_iarg_43_din1),
        .ap_bram_43_dout1(ap_bram_iarg_43_dout1),
        .ap_bram_43_we1(ap_bram_iarg_43_we1),
        .ap_bram_43_en1(ap_bram_iarg_43_en1),
        .s_axis_bram_44_tlast(s_axis_bram_44_tlast),
        .s_axis_bram_44_tvalid(s_axis_bram_44_tvalid),
        .s_axis_bram_44_tkeep(s_axis_bram_44_tkeep),
        .s_axis_bram_44_tstrb(s_axis_bram_44_tstrb),
        .s_axis_bram_44_tdata(s_axis_bram_44_tdata),
        .s_axis_bram_44_tready(s_axis_bram_44_tready),
        .ap_bram_44_addr0(ap_bram_iarg_44_addr0),
        .ap_bram_44_din0(ap_bram_iarg_44_din0),
        .ap_bram_44_dout0(ap_bram_iarg_44_dout0),
        .ap_bram_44_we0(ap_bram_iarg_44_we0),
        .ap_bram_44_en0(ap_bram_iarg_44_en0),
        .ap_bram_44_addr1(ap_bram_iarg_44_addr1),
        .ap_bram_44_din1(ap_bram_iarg_44_din1),
        .ap_bram_44_dout1(ap_bram_iarg_44_dout1),
        .ap_bram_44_we1(ap_bram_iarg_44_we1),
        .ap_bram_44_en1(ap_bram_iarg_44_en1),
        .s_axis_bram_45_tlast(s_axis_bram_45_tlast),
        .s_axis_bram_45_tvalid(s_axis_bram_45_tvalid),
        .s_axis_bram_45_tkeep(s_axis_bram_45_tkeep),
        .s_axis_bram_45_tstrb(s_axis_bram_45_tstrb),
        .s_axis_bram_45_tdata(s_axis_bram_45_tdata),
        .s_axis_bram_45_tready(s_axis_bram_45_tready),
        .ap_bram_45_addr0(ap_bram_iarg_45_addr0),
        .ap_bram_45_din0(ap_bram_iarg_45_din0),
        .ap_bram_45_dout0(ap_bram_iarg_45_dout0),
        .ap_bram_45_we0(ap_bram_iarg_45_we0),
        .ap_bram_45_en0(ap_bram_iarg_45_en0),
        .ap_bram_45_addr1(ap_bram_iarg_45_addr1),
        .ap_bram_45_din1(ap_bram_iarg_45_din1),
        .ap_bram_45_dout1(ap_bram_iarg_45_dout1),
        .ap_bram_45_we1(ap_bram_iarg_45_we1),
        .ap_bram_45_en1(ap_bram_iarg_45_en1),
        .s_axis_bram_46_tlast(s_axis_bram_46_tlast),
        .s_axis_bram_46_tvalid(s_axis_bram_46_tvalid),
        .s_axis_bram_46_tkeep(s_axis_bram_46_tkeep),
        .s_axis_bram_46_tstrb(s_axis_bram_46_tstrb),
        .s_axis_bram_46_tdata(s_axis_bram_46_tdata),
        .s_axis_bram_46_tready(s_axis_bram_46_tready),
        .ap_bram_46_addr0(ap_bram_iarg_46_addr0),
        .ap_bram_46_din0(ap_bram_iarg_46_din0),
        .ap_bram_46_dout0(ap_bram_iarg_46_dout0),
        .ap_bram_46_we0(ap_bram_iarg_46_we0),
        .ap_bram_46_en0(ap_bram_iarg_46_en0),
        .ap_bram_46_addr1(ap_bram_iarg_46_addr1),
        .ap_bram_46_din1(ap_bram_iarg_46_din1),
        .ap_bram_46_dout1(ap_bram_iarg_46_dout1),
        .ap_bram_46_we1(ap_bram_iarg_46_we1),
        .ap_bram_46_en1(ap_bram_iarg_46_en1),
        .s_axis_bram_47_tlast(s_axis_bram_47_tlast),
        .s_axis_bram_47_tvalid(s_axis_bram_47_tvalid),
        .s_axis_bram_47_tkeep(s_axis_bram_47_tkeep),
        .s_axis_bram_47_tstrb(s_axis_bram_47_tstrb),
        .s_axis_bram_47_tdata(s_axis_bram_47_tdata),
        .s_axis_bram_47_tready(s_axis_bram_47_tready),
        .ap_bram_47_addr0(ap_bram_iarg_47_addr0),
        .ap_bram_47_din0(ap_bram_iarg_47_din0),
        .ap_bram_47_dout0(ap_bram_iarg_47_dout0),
        .ap_bram_47_we0(ap_bram_iarg_47_we0),
        .ap_bram_47_en0(ap_bram_iarg_47_en0),
        .ap_bram_47_addr1(ap_bram_iarg_47_addr1),
        .ap_bram_47_din1(ap_bram_iarg_47_din1),
        .ap_bram_47_dout1(ap_bram_iarg_47_dout1),
        .ap_bram_47_we1(ap_bram_iarg_47_we1),
        .ap_bram_47_en1(ap_bram_iarg_47_en1),
        .s_axis_bram_48_tlast(s_axis_bram_48_tlast),
        .s_axis_bram_48_tvalid(s_axis_bram_48_tvalid),
        .s_axis_bram_48_tkeep(s_axis_bram_48_tkeep),
        .s_axis_bram_48_tstrb(s_axis_bram_48_tstrb),
        .s_axis_bram_48_tdata(s_axis_bram_48_tdata),
        .s_axis_bram_48_tready(s_axis_bram_48_tready),
        .ap_bram_48_addr0(ap_bram_iarg_48_addr0),
        .ap_bram_48_din0(ap_bram_iarg_48_din0),
        .ap_bram_48_dout0(ap_bram_iarg_48_dout0),
        .ap_bram_48_we0(ap_bram_iarg_48_we0),
        .ap_bram_48_en0(ap_bram_iarg_48_en0),
        .ap_bram_48_addr1(ap_bram_iarg_48_addr1),
        .ap_bram_48_din1(ap_bram_iarg_48_din1),
        .ap_bram_48_dout1(ap_bram_iarg_48_dout1),
        .ap_bram_48_we1(ap_bram_iarg_48_we1),
        .ap_bram_48_en1(ap_bram_iarg_48_en1),
        .s_axis_bram_49_tlast(s_axis_bram_49_tlast),
        .s_axis_bram_49_tvalid(s_axis_bram_49_tvalid),
        .s_axis_bram_49_tkeep(s_axis_bram_49_tkeep),
        .s_axis_bram_49_tstrb(s_axis_bram_49_tstrb),
        .s_axis_bram_49_tdata(s_axis_bram_49_tdata),
        .s_axis_bram_49_tready(s_axis_bram_49_tready),
        .ap_bram_49_addr0(ap_bram_iarg_49_addr0),
        .ap_bram_49_din0(ap_bram_iarg_49_din0),
        .ap_bram_49_dout0(ap_bram_iarg_49_dout0),
        .ap_bram_49_we0(ap_bram_iarg_49_we0),
        .ap_bram_49_en0(ap_bram_iarg_49_en0),
        .ap_bram_49_addr1(ap_bram_iarg_49_addr1),
        .ap_bram_49_din1(ap_bram_iarg_49_din1),
        .ap_bram_49_dout1(ap_bram_iarg_49_dout1),
        .ap_bram_49_we1(ap_bram_iarg_49_we1),
        .ap_bram_49_en1(ap_bram_iarg_49_en1),
        .s_axis_bram_50_tlast(s_axis_bram_50_tlast),
        .s_axis_bram_50_tvalid(s_axis_bram_50_tvalid),
        .s_axis_bram_50_tkeep(s_axis_bram_50_tkeep),
        .s_axis_bram_50_tstrb(s_axis_bram_50_tstrb),
        .s_axis_bram_50_tdata(s_axis_bram_50_tdata),
        .s_axis_bram_50_tready(s_axis_bram_50_tready),
        .ap_bram_50_addr0(ap_bram_iarg_50_addr0),
        .ap_bram_50_din0(ap_bram_iarg_50_din0),
        .ap_bram_50_dout0(ap_bram_iarg_50_dout0),
        .ap_bram_50_we0(ap_bram_iarg_50_we0),
        .ap_bram_50_en0(ap_bram_iarg_50_en0),
        .ap_bram_50_addr1(ap_bram_iarg_50_addr1),
        .ap_bram_50_din1(ap_bram_iarg_50_din1),
        .ap_bram_50_dout1(ap_bram_iarg_50_dout1),
        .ap_bram_50_we1(ap_bram_iarg_50_we1),
        .ap_bram_50_en1(ap_bram_iarg_50_en1),
        .s_axis_bram_51_tlast(s_axis_bram_51_tlast),
        .s_axis_bram_51_tvalid(s_axis_bram_51_tvalid),
        .s_axis_bram_51_tkeep(s_axis_bram_51_tkeep),
        .s_axis_bram_51_tstrb(s_axis_bram_51_tstrb),
        .s_axis_bram_51_tdata(s_axis_bram_51_tdata),
        .s_axis_bram_51_tready(s_axis_bram_51_tready),
        .ap_bram_51_addr0(ap_bram_iarg_51_addr0),
        .ap_bram_51_din0(ap_bram_iarg_51_din0),
        .ap_bram_51_dout0(ap_bram_iarg_51_dout0),
        .ap_bram_51_we0(ap_bram_iarg_51_we0),
        .ap_bram_51_en0(ap_bram_iarg_51_en0),
        .ap_bram_51_addr1(ap_bram_iarg_51_addr1),
        .ap_bram_51_din1(ap_bram_iarg_51_din1),
        .ap_bram_51_dout1(ap_bram_iarg_51_dout1),
        .ap_bram_51_we1(ap_bram_iarg_51_we1),
        .ap_bram_51_en1(ap_bram_iarg_51_en1),
        .s_axis_bram_52_tlast(s_axis_bram_52_tlast),
        .s_axis_bram_52_tvalid(s_axis_bram_52_tvalid),
        .s_axis_bram_52_tkeep(s_axis_bram_52_tkeep),
        .s_axis_bram_52_tstrb(s_axis_bram_52_tstrb),
        .s_axis_bram_52_tdata(s_axis_bram_52_tdata),
        .s_axis_bram_52_tready(s_axis_bram_52_tready),
        .ap_bram_52_addr0(ap_bram_iarg_52_addr0),
        .ap_bram_52_din0(ap_bram_iarg_52_din0),
        .ap_bram_52_dout0(ap_bram_iarg_52_dout0),
        .ap_bram_52_we0(ap_bram_iarg_52_we0),
        .ap_bram_52_en0(ap_bram_iarg_52_en0),
        .ap_bram_52_addr1(ap_bram_iarg_52_addr1),
        .ap_bram_52_din1(ap_bram_iarg_52_din1),
        .ap_bram_52_dout1(ap_bram_iarg_52_dout1),
        .ap_bram_52_we1(ap_bram_iarg_52_we1),
        .ap_bram_52_en1(ap_bram_iarg_52_en1),
        .s_axis_bram_53_tlast(s_axis_bram_53_tlast),
        .s_axis_bram_53_tvalid(s_axis_bram_53_tvalid),
        .s_axis_bram_53_tkeep(s_axis_bram_53_tkeep),
        .s_axis_bram_53_tstrb(s_axis_bram_53_tstrb),
        .s_axis_bram_53_tdata(s_axis_bram_53_tdata),
        .s_axis_bram_53_tready(s_axis_bram_53_tready),
        .ap_bram_53_addr0(ap_bram_iarg_53_addr0),
        .ap_bram_53_din0(ap_bram_iarg_53_din0),
        .ap_bram_53_dout0(ap_bram_iarg_53_dout0),
        .ap_bram_53_we0(ap_bram_iarg_53_we0),
        .ap_bram_53_en0(ap_bram_iarg_53_en0),
        .ap_bram_53_addr1(ap_bram_iarg_53_addr1),
        .ap_bram_53_din1(ap_bram_iarg_53_din1),
        .ap_bram_53_dout1(ap_bram_iarg_53_dout1),
        .ap_bram_53_we1(ap_bram_iarg_53_we1),
        .ap_bram_53_en1(ap_bram_iarg_53_en1),
        .s_axis_bram_54_tlast(s_axis_bram_54_tlast),
        .s_axis_bram_54_tvalid(s_axis_bram_54_tvalid),
        .s_axis_bram_54_tkeep(s_axis_bram_54_tkeep),
        .s_axis_bram_54_tstrb(s_axis_bram_54_tstrb),
        .s_axis_bram_54_tdata(s_axis_bram_54_tdata),
        .s_axis_bram_54_tready(s_axis_bram_54_tready),
        .ap_bram_54_addr0(ap_bram_iarg_54_addr0),
        .ap_bram_54_din0(ap_bram_iarg_54_din0),
        .ap_bram_54_dout0(ap_bram_iarg_54_dout0),
        .ap_bram_54_we0(ap_bram_iarg_54_we0),
        .ap_bram_54_en0(ap_bram_iarg_54_en0),
        .ap_bram_54_addr1(ap_bram_iarg_54_addr1),
        .ap_bram_54_din1(ap_bram_iarg_54_din1),
        .ap_bram_54_dout1(ap_bram_iarg_54_dout1),
        .ap_bram_54_we1(ap_bram_iarg_54_we1),
        .ap_bram_54_en1(ap_bram_iarg_54_en1),
        .s_axis_bram_55_tlast(s_axis_bram_55_tlast),
        .s_axis_bram_55_tvalid(s_axis_bram_55_tvalid),
        .s_axis_bram_55_tkeep(s_axis_bram_55_tkeep),
        .s_axis_bram_55_tstrb(s_axis_bram_55_tstrb),
        .s_axis_bram_55_tdata(s_axis_bram_55_tdata),
        .s_axis_bram_55_tready(s_axis_bram_55_tready),
        .ap_bram_55_addr0(ap_bram_iarg_55_addr0),
        .ap_bram_55_din0(ap_bram_iarg_55_din0),
        .ap_bram_55_dout0(ap_bram_iarg_55_dout0),
        .ap_bram_55_we0(ap_bram_iarg_55_we0),
        .ap_bram_55_en0(ap_bram_iarg_55_en0),
        .ap_bram_55_addr1(ap_bram_iarg_55_addr1),
        .ap_bram_55_din1(ap_bram_iarg_55_din1),
        .ap_bram_55_dout1(ap_bram_iarg_55_dout1),
        .ap_bram_55_we1(ap_bram_iarg_55_we1),
        .ap_bram_55_en1(ap_bram_iarg_55_en1),
        .s_axis_bram_56_tlast(s_axis_bram_56_tlast),
        .s_axis_bram_56_tvalid(s_axis_bram_56_tvalid),
        .s_axis_bram_56_tkeep(s_axis_bram_56_tkeep),
        .s_axis_bram_56_tstrb(s_axis_bram_56_tstrb),
        .s_axis_bram_56_tdata(s_axis_bram_56_tdata),
        .s_axis_bram_56_tready(s_axis_bram_56_tready),
        .ap_bram_56_addr0(ap_bram_iarg_56_addr0),
        .ap_bram_56_din0(ap_bram_iarg_56_din0),
        .ap_bram_56_dout0(ap_bram_iarg_56_dout0),
        .ap_bram_56_we0(ap_bram_iarg_56_we0),
        .ap_bram_56_en0(ap_bram_iarg_56_en0),
        .ap_bram_56_addr1(ap_bram_iarg_56_addr1),
        .ap_bram_56_din1(ap_bram_iarg_56_din1),
        .ap_bram_56_dout1(ap_bram_iarg_56_dout1),
        .ap_bram_56_we1(ap_bram_iarg_56_we1),
        .ap_bram_56_en1(ap_bram_iarg_56_en1),
        .s_axis_bram_57_tlast(s_axis_bram_57_tlast),
        .s_axis_bram_57_tvalid(s_axis_bram_57_tvalid),
        .s_axis_bram_57_tkeep(s_axis_bram_57_tkeep),
        .s_axis_bram_57_tstrb(s_axis_bram_57_tstrb),
        .s_axis_bram_57_tdata(s_axis_bram_57_tdata),
        .s_axis_bram_57_tready(s_axis_bram_57_tready),
        .ap_bram_57_addr0(ap_bram_iarg_57_addr0),
        .ap_bram_57_din0(ap_bram_iarg_57_din0),
        .ap_bram_57_dout0(ap_bram_iarg_57_dout0),
        .ap_bram_57_we0(ap_bram_iarg_57_we0),
        .ap_bram_57_en0(ap_bram_iarg_57_en0),
        .ap_bram_57_addr1(ap_bram_iarg_57_addr1),
        .ap_bram_57_din1(ap_bram_iarg_57_din1),
        .ap_bram_57_dout1(ap_bram_iarg_57_dout1),
        .ap_bram_57_we1(ap_bram_iarg_57_we1),
        .ap_bram_57_en1(ap_bram_iarg_57_en1),
        .s_axis_bram_58_tlast(s_axis_bram_58_tlast),
        .s_axis_bram_58_tvalid(s_axis_bram_58_tvalid),
        .s_axis_bram_58_tkeep(s_axis_bram_58_tkeep),
        .s_axis_bram_58_tstrb(s_axis_bram_58_tstrb),
        .s_axis_bram_58_tdata(s_axis_bram_58_tdata),
        .s_axis_bram_58_tready(s_axis_bram_58_tready),
        .ap_bram_58_addr0(ap_bram_iarg_58_addr0),
        .ap_bram_58_din0(ap_bram_iarg_58_din0),
        .ap_bram_58_dout0(ap_bram_iarg_58_dout0),
        .ap_bram_58_we0(ap_bram_iarg_58_we0),
        .ap_bram_58_en0(ap_bram_iarg_58_en0),
        .ap_bram_58_addr1(ap_bram_iarg_58_addr1),
        .ap_bram_58_din1(ap_bram_iarg_58_din1),
        .ap_bram_58_dout1(ap_bram_iarg_58_dout1),
        .ap_bram_58_we1(ap_bram_iarg_58_we1),
        .ap_bram_58_en1(ap_bram_iarg_58_en1),
        .s_axis_bram_59_tlast(s_axis_bram_59_tlast),
        .s_axis_bram_59_tvalid(s_axis_bram_59_tvalid),
        .s_axis_bram_59_tkeep(s_axis_bram_59_tkeep),
        .s_axis_bram_59_tstrb(s_axis_bram_59_tstrb),
        .s_axis_bram_59_tdata(s_axis_bram_59_tdata),
        .s_axis_bram_59_tready(s_axis_bram_59_tready),
        .ap_bram_59_addr0(ap_bram_iarg_59_addr0),
        .ap_bram_59_din0(ap_bram_iarg_59_din0),
        .ap_bram_59_dout0(ap_bram_iarg_59_dout0),
        .ap_bram_59_we0(ap_bram_iarg_59_we0),
        .ap_bram_59_en0(ap_bram_iarg_59_en0),
        .ap_bram_59_addr1(ap_bram_iarg_59_addr1),
        .ap_bram_59_din1(ap_bram_iarg_59_din1),
        .ap_bram_59_dout1(ap_bram_iarg_59_dout1),
        .ap_bram_59_we1(ap_bram_iarg_59_we1),
        .ap_bram_59_en1(ap_bram_iarg_59_en1),
        .s_axis_bram_60_tlast(s_axis_bram_60_tlast),
        .s_axis_bram_60_tvalid(s_axis_bram_60_tvalid),
        .s_axis_bram_60_tkeep(s_axis_bram_60_tkeep),
        .s_axis_bram_60_tstrb(s_axis_bram_60_tstrb),
        .s_axis_bram_60_tdata(s_axis_bram_60_tdata),
        .s_axis_bram_60_tready(s_axis_bram_60_tready),
        .ap_bram_60_addr0(ap_bram_iarg_60_addr0),
        .ap_bram_60_din0(ap_bram_iarg_60_din0),
        .ap_bram_60_dout0(ap_bram_iarg_60_dout0),
        .ap_bram_60_we0(ap_bram_iarg_60_we0),
        .ap_bram_60_en0(ap_bram_iarg_60_en0),
        .ap_bram_60_addr1(ap_bram_iarg_60_addr1),
        .ap_bram_60_din1(ap_bram_iarg_60_din1),
        .ap_bram_60_dout1(ap_bram_iarg_60_dout1),
        .ap_bram_60_we1(ap_bram_iarg_60_we1),
        .ap_bram_60_en1(ap_bram_iarg_60_en1),
        .s_axis_bram_61_tlast(s_axis_bram_61_tlast),
        .s_axis_bram_61_tvalid(s_axis_bram_61_tvalid),
        .s_axis_bram_61_tkeep(s_axis_bram_61_tkeep),
        .s_axis_bram_61_tstrb(s_axis_bram_61_tstrb),
        .s_axis_bram_61_tdata(s_axis_bram_61_tdata),
        .s_axis_bram_61_tready(s_axis_bram_61_tready),
        .ap_bram_61_addr0(ap_bram_iarg_61_addr0),
        .ap_bram_61_din0(ap_bram_iarg_61_din0),
        .ap_bram_61_dout0(ap_bram_iarg_61_dout0),
        .ap_bram_61_we0(ap_bram_iarg_61_we0),
        .ap_bram_61_en0(ap_bram_iarg_61_en0),
        .ap_bram_61_addr1(ap_bram_iarg_61_addr1),
        .ap_bram_61_din1(ap_bram_iarg_61_din1),
        .ap_bram_61_dout1(ap_bram_iarg_61_dout1),
        .ap_bram_61_we1(ap_bram_iarg_61_we1),
        .ap_bram_61_en1(ap_bram_iarg_61_en1),
        .s_axis_bram_62_tlast(s_axis_bram_62_tlast),
        .s_axis_bram_62_tvalid(s_axis_bram_62_tvalid),
        .s_axis_bram_62_tkeep(s_axis_bram_62_tkeep),
        .s_axis_bram_62_tstrb(s_axis_bram_62_tstrb),
        .s_axis_bram_62_tdata(s_axis_bram_62_tdata),
        .s_axis_bram_62_tready(s_axis_bram_62_tready),
        .ap_bram_62_addr0(ap_bram_iarg_62_addr0),
        .ap_bram_62_din0(ap_bram_iarg_62_din0),
        .ap_bram_62_dout0(ap_bram_iarg_62_dout0),
        .ap_bram_62_we0(ap_bram_iarg_62_we0),
        .ap_bram_62_en0(ap_bram_iarg_62_en0),
        .ap_bram_62_addr1(ap_bram_iarg_62_addr1),
        .ap_bram_62_din1(ap_bram_iarg_62_din1),
        .ap_bram_62_dout1(ap_bram_iarg_62_dout1),
        .ap_bram_62_we1(ap_bram_iarg_62_we1),
        .ap_bram_62_en1(ap_bram_iarg_62_en1),
        .s_axis_bram_63_tlast(s_axis_bram_63_tlast),
        .s_axis_bram_63_tvalid(s_axis_bram_63_tvalid),
        .s_axis_bram_63_tkeep(s_axis_bram_63_tkeep),
        .s_axis_bram_63_tstrb(s_axis_bram_63_tstrb),
        .s_axis_bram_63_tdata(s_axis_bram_63_tdata),
        .s_axis_bram_63_tready(s_axis_bram_63_tready),
        .ap_bram_63_addr0(ap_bram_iarg_63_addr0),
        .ap_bram_63_din0(ap_bram_iarg_63_din0),
        .ap_bram_63_dout0(ap_bram_iarg_63_dout0),
        .ap_bram_63_we0(ap_bram_iarg_63_we0),
        .ap_bram_63_en0(ap_bram_iarg_63_en0),
        .ap_bram_63_addr1(ap_bram_iarg_63_addr1),
        .ap_bram_63_din1(ap_bram_iarg_63_din1),
        .ap_bram_63_dout1(ap_bram_iarg_63_dout1),
        .ap_bram_63_we1(ap_bram_iarg_63_we1),
        .ap_bram_63_en1(ap_bram_iarg_63_en1),
        .s_axis_bram_64_tlast(s_axis_bram_64_tlast),
        .s_axis_bram_64_tvalid(s_axis_bram_64_tvalid),
        .s_axis_bram_64_tkeep(s_axis_bram_64_tkeep),
        .s_axis_bram_64_tstrb(s_axis_bram_64_tstrb),
        .s_axis_bram_64_tdata(s_axis_bram_64_tdata),
        .s_axis_bram_64_tready(s_axis_bram_64_tready),
        .ap_bram_64_addr0(ap_bram_iarg_64_addr0),
        .ap_bram_64_din0(ap_bram_iarg_64_din0),
        .ap_bram_64_dout0(ap_bram_iarg_64_dout0),
        .ap_bram_64_we0(ap_bram_iarg_64_we0),
        .ap_bram_64_en0(ap_bram_iarg_64_en0),
        .ap_bram_64_addr1(ap_bram_iarg_64_addr1),
        .ap_bram_64_din1(ap_bram_iarg_64_din1),
        .ap_bram_64_dout1(ap_bram_iarg_64_dout1),
        .ap_bram_64_we1(ap_bram_iarg_64_we1),
        .ap_bram_64_en1(ap_bram_iarg_64_en1),
        .s_axis_bram_65_tlast(s_axis_bram_65_tlast),
        .s_axis_bram_65_tvalid(s_axis_bram_65_tvalid),
        .s_axis_bram_65_tkeep(s_axis_bram_65_tkeep),
        .s_axis_bram_65_tstrb(s_axis_bram_65_tstrb),
        .s_axis_bram_65_tdata(s_axis_bram_65_tdata),
        .s_axis_bram_65_tready(s_axis_bram_65_tready),
        .ap_bram_65_addr0(ap_bram_iarg_65_addr0),
        .ap_bram_65_din0(ap_bram_iarg_65_din0),
        .ap_bram_65_dout0(ap_bram_iarg_65_dout0),
        .ap_bram_65_we0(ap_bram_iarg_65_we0),
        .ap_bram_65_en0(ap_bram_iarg_65_en0),
        .ap_bram_65_addr1(ap_bram_iarg_65_addr1),
        .ap_bram_65_din1(ap_bram_iarg_65_din1),
        .ap_bram_65_dout1(ap_bram_iarg_65_dout1),
        .ap_bram_65_we1(ap_bram_iarg_65_we1),
        .ap_bram_65_en1(ap_bram_iarg_65_en1),
        .s_axis_bram_66_tlast(s_axis_bram_66_tlast),
        .s_axis_bram_66_tvalid(s_axis_bram_66_tvalid),
        .s_axis_bram_66_tkeep(s_axis_bram_66_tkeep),
        .s_axis_bram_66_tstrb(s_axis_bram_66_tstrb),
        .s_axis_bram_66_tdata(s_axis_bram_66_tdata),
        .s_axis_bram_66_tready(s_axis_bram_66_tready),
        .ap_bram_66_addr0(ap_bram_iarg_66_addr0),
        .ap_bram_66_din0(ap_bram_iarg_66_din0),
        .ap_bram_66_dout0(ap_bram_iarg_66_dout0),
        .ap_bram_66_we0(ap_bram_iarg_66_we0),
        .ap_bram_66_en0(ap_bram_iarg_66_en0),
        .ap_bram_66_addr1(ap_bram_iarg_66_addr1),
        .ap_bram_66_din1(ap_bram_iarg_66_din1),
        .ap_bram_66_dout1(ap_bram_iarg_66_dout1),
        .ap_bram_66_we1(ap_bram_iarg_66_we1),
        .ap_bram_66_en1(ap_bram_iarg_66_en1),
        .s_axis_bram_67_tlast(s_axis_bram_67_tlast),
        .s_axis_bram_67_tvalid(s_axis_bram_67_tvalid),
        .s_axis_bram_67_tkeep(s_axis_bram_67_tkeep),
        .s_axis_bram_67_tstrb(s_axis_bram_67_tstrb),
        .s_axis_bram_67_tdata(s_axis_bram_67_tdata),
        .s_axis_bram_67_tready(s_axis_bram_67_tready),
        .ap_bram_67_addr0(ap_bram_iarg_67_addr0),
        .ap_bram_67_din0(ap_bram_iarg_67_din0),
        .ap_bram_67_dout0(ap_bram_iarg_67_dout0),
        .ap_bram_67_we0(ap_bram_iarg_67_we0),
        .ap_bram_67_en0(ap_bram_iarg_67_en0),
        .ap_bram_67_addr1(ap_bram_iarg_67_addr1),
        .ap_bram_67_din1(ap_bram_iarg_67_din1),
        .ap_bram_67_dout1(ap_bram_iarg_67_dout1),
        .ap_bram_67_we1(ap_bram_iarg_67_we1),
        .ap_bram_67_en1(ap_bram_iarg_67_en1),
        .s_axis_bram_68_tlast(s_axis_bram_68_tlast),
        .s_axis_bram_68_tvalid(s_axis_bram_68_tvalid),
        .s_axis_bram_68_tkeep(s_axis_bram_68_tkeep),
        .s_axis_bram_68_tstrb(s_axis_bram_68_tstrb),
        .s_axis_bram_68_tdata(s_axis_bram_68_tdata),
        .s_axis_bram_68_tready(s_axis_bram_68_tready),
        .ap_bram_68_addr0(ap_bram_iarg_68_addr0),
        .ap_bram_68_din0(ap_bram_iarg_68_din0),
        .ap_bram_68_dout0(ap_bram_iarg_68_dout0),
        .ap_bram_68_we0(ap_bram_iarg_68_we0),
        .ap_bram_68_en0(ap_bram_iarg_68_en0),
        .ap_bram_68_addr1(ap_bram_iarg_68_addr1),
        .ap_bram_68_din1(ap_bram_iarg_68_din1),
        .ap_bram_68_dout1(ap_bram_iarg_68_dout1),
        .ap_bram_68_we1(ap_bram_iarg_68_we1),
        .ap_bram_68_en1(ap_bram_iarg_68_en1),
        .s_axis_bram_69_tlast(s_axis_bram_69_tlast),
        .s_axis_bram_69_tvalid(s_axis_bram_69_tvalid),
        .s_axis_bram_69_tkeep(s_axis_bram_69_tkeep),
        .s_axis_bram_69_tstrb(s_axis_bram_69_tstrb),
        .s_axis_bram_69_tdata(s_axis_bram_69_tdata),
        .s_axis_bram_69_tready(s_axis_bram_69_tready),
        .ap_bram_69_addr0(ap_bram_iarg_69_addr0),
        .ap_bram_69_din0(ap_bram_iarg_69_din0),
        .ap_bram_69_dout0(ap_bram_iarg_69_dout0),
        .ap_bram_69_we0(ap_bram_iarg_69_we0),
        .ap_bram_69_en0(ap_bram_iarg_69_en0),
        .ap_bram_69_addr1(ap_bram_iarg_69_addr1),
        .ap_bram_69_din1(ap_bram_iarg_69_din1),
        .ap_bram_69_dout1(ap_bram_iarg_69_dout1),
        .ap_bram_69_we1(ap_bram_iarg_69_we1),
        .ap_bram_69_en1(ap_bram_iarg_69_en1),
        .s_axis_bram_70_tlast(s_axis_bram_70_tlast),
        .s_axis_bram_70_tvalid(s_axis_bram_70_tvalid),
        .s_axis_bram_70_tkeep(s_axis_bram_70_tkeep),
        .s_axis_bram_70_tstrb(s_axis_bram_70_tstrb),
        .s_axis_bram_70_tdata(s_axis_bram_70_tdata),
        .s_axis_bram_70_tready(s_axis_bram_70_tready),
        .ap_bram_70_addr0(ap_bram_iarg_70_addr0),
        .ap_bram_70_din0(ap_bram_iarg_70_din0),
        .ap_bram_70_dout0(ap_bram_iarg_70_dout0),
        .ap_bram_70_we0(ap_bram_iarg_70_we0),
        .ap_bram_70_en0(ap_bram_iarg_70_en0),
        .ap_bram_70_addr1(ap_bram_iarg_70_addr1),
        .ap_bram_70_din1(ap_bram_iarg_70_din1),
        .ap_bram_70_dout1(ap_bram_iarg_70_dout1),
        .ap_bram_70_we1(ap_bram_iarg_70_we1),
        .ap_bram_70_en1(ap_bram_iarg_70_en1),
        .s_axis_bram_71_tlast(s_axis_bram_71_tlast),
        .s_axis_bram_71_tvalid(s_axis_bram_71_tvalid),
        .s_axis_bram_71_tkeep(s_axis_bram_71_tkeep),
        .s_axis_bram_71_tstrb(s_axis_bram_71_tstrb),
        .s_axis_bram_71_tdata(s_axis_bram_71_tdata),
        .s_axis_bram_71_tready(s_axis_bram_71_tready),
        .ap_bram_71_addr0(ap_bram_iarg_71_addr0),
        .ap_bram_71_din0(ap_bram_iarg_71_din0),
        .ap_bram_71_dout0(ap_bram_iarg_71_dout0),
        .ap_bram_71_we0(ap_bram_iarg_71_we0),
        .ap_bram_71_en0(ap_bram_iarg_71_en0),
        .ap_bram_71_addr1(ap_bram_iarg_71_addr1),
        .ap_bram_71_din1(ap_bram_iarg_71_din1),
        .ap_bram_71_dout1(ap_bram_iarg_71_dout1),
        .ap_bram_71_we1(ap_bram_iarg_71_we1),
        .ap_bram_71_en1(ap_bram_iarg_71_en1),
        .s_axis_bram_72_tlast(s_axis_bram_72_tlast),
        .s_axis_bram_72_tvalid(s_axis_bram_72_tvalid),
        .s_axis_bram_72_tkeep(s_axis_bram_72_tkeep),
        .s_axis_bram_72_tstrb(s_axis_bram_72_tstrb),
        .s_axis_bram_72_tdata(s_axis_bram_72_tdata),
        .s_axis_bram_72_tready(s_axis_bram_72_tready),
        .ap_bram_72_addr0(ap_bram_iarg_72_addr0),
        .ap_bram_72_din0(ap_bram_iarg_72_din0),
        .ap_bram_72_dout0(ap_bram_iarg_72_dout0),
        .ap_bram_72_we0(ap_bram_iarg_72_we0),
        .ap_bram_72_en0(ap_bram_iarg_72_en0),
        .ap_bram_72_addr1(ap_bram_iarg_72_addr1),
        .ap_bram_72_din1(ap_bram_iarg_72_din1),
        .ap_bram_72_dout1(ap_bram_iarg_72_dout1),
        .ap_bram_72_we1(ap_bram_iarg_72_we1),
        .ap_bram_72_en1(ap_bram_iarg_72_en1),
        .s_axis_bram_73_tlast(s_axis_bram_73_tlast),
        .s_axis_bram_73_tvalid(s_axis_bram_73_tvalid),
        .s_axis_bram_73_tkeep(s_axis_bram_73_tkeep),
        .s_axis_bram_73_tstrb(s_axis_bram_73_tstrb),
        .s_axis_bram_73_tdata(s_axis_bram_73_tdata),
        .s_axis_bram_73_tready(s_axis_bram_73_tready),
        .ap_bram_73_addr0(ap_bram_iarg_73_addr0),
        .ap_bram_73_din0(ap_bram_iarg_73_din0),
        .ap_bram_73_dout0(ap_bram_iarg_73_dout0),
        .ap_bram_73_we0(ap_bram_iarg_73_we0),
        .ap_bram_73_en0(ap_bram_iarg_73_en0),
        .ap_bram_73_addr1(ap_bram_iarg_73_addr1),
        .ap_bram_73_din1(ap_bram_iarg_73_din1),
        .ap_bram_73_dout1(ap_bram_iarg_73_dout1),
        .ap_bram_73_we1(ap_bram_iarg_73_we1),
        .ap_bram_73_en1(ap_bram_iarg_73_en1),
        .s_axis_bram_74_tlast(s_axis_bram_74_tlast),
        .s_axis_bram_74_tvalid(s_axis_bram_74_tvalid),
        .s_axis_bram_74_tkeep(s_axis_bram_74_tkeep),
        .s_axis_bram_74_tstrb(s_axis_bram_74_tstrb),
        .s_axis_bram_74_tdata(s_axis_bram_74_tdata),
        .s_axis_bram_74_tready(s_axis_bram_74_tready),
        .ap_bram_74_addr0(ap_bram_iarg_74_addr0),
        .ap_bram_74_din0(ap_bram_iarg_74_din0),
        .ap_bram_74_dout0(ap_bram_iarg_74_dout0),
        .ap_bram_74_we0(ap_bram_iarg_74_we0),
        .ap_bram_74_en0(ap_bram_iarg_74_en0),
        .ap_bram_74_addr1(ap_bram_iarg_74_addr1),
        .ap_bram_74_din1(ap_bram_iarg_74_din1),
        .ap_bram_74_dout1(ap_bram_iarg_74_dout1),
        .ap_bram_74_we1(ap_bram_iarg_74_we1),
        .ap_bram_74_en1(ap_bram_iarg_74_en1),
        .s_axis_bram_75_tlast(s_axis_bram_75_tlast),
        .s_axis_bram_75_tvalid(s_axis_bram_75_tvalid),
        .s_axis_bram_75_tkeep(s_axis_bram_75_tkeep),
        .s_axis_bram_75_tstrb(s_axis_bram_75_tstrb),
        .s_axis_bram_75_tdata(s_axis_bram_75_tdata),
        .s_axis_bram_75_tready(s_axis_bram_75_tready),
        .ap_bram_75_addr0(ap_bram_iarg_75_addr0),
        .ap_bram_75_din0(ap_bram_iarg_75_din0),
        .ap_bram_75_dout0(ap_bram_iarg_75_dout0),
        .ap_bram_75_we0(ap_bram_iarg_75_we0),
        .ap_bram_75_en0(ap_bram_iarg_75_en0),
        .ap_bram_75_addr1(ap_bram_iarg_75_addr1),
        .ap_bram_75_din1(ap_bram_iarg_75_din1),
        .ap_bram_75_dout1(ap_bram_iarg_75_dout1),
        .ap_bram_75_we1(ap_bram_iarg_75_we1),
        .ap_bram_75_en1(ap_bram_iarg_75_en1),
        .s_axis_bram_76_tlast(s_axis_bram_76_tlast),
        .s_axis_bram_76_tvalid(s_axis_bram_76_tvalid),
        .s_axis_bram_76_tkeep(s_axis_bram_76_tkeep),
        .s_axis_bram_76_tstrb(s_axis_bram_76_tstrb),
        .s_axis_bram_76_tdata(s_axis_bram_76_tdata),
        .s_axis_bram_76_tready(s_axis_bram_76_tready),
        .ap_bram_76_addr0(ap_bram_iarg_76_addr0),
        .ap_bram_76_din0(ap_bram_iarg_76_din0),
        .ap_bram_76_dout0(ap_bram_iarg_76_dout0),
        .ap_bram_76_we0(ap_bram_iarg_76_we0),
        .ap_bram_76_en0(ap_bram_iarg_76_en0),
        .ap_bram_76_addr1(ap_bram_iarg_76_addr1),
        .ap_bram_76_din1(ap_bram_iarg_76_din1),
        .ap_bram_76_dout1(ap_bram_iarg_76_dout1),
        .ap_bram_76_we1(ap_bram_iarg_76_we1),
        .ap_bram_76_en1(ap_bram_iarg_76_en1),
        .s_axis_bram_77_tlast(s_axis_bram_77_tlast),
        .s_axis_bram_77_tvalid(s_axis_bram_77_tvalid),
        .s_axis_bram_77_tkeep(s_axis_bram_77_tkeep),
        .s_axis_bram_77_tstrb(s_axis_bram_77_tstrb),
        .s_axis_bram_77_tdata(s_axis_bram_77_tdata),
        .s_axis_bram_77_tready(s_axis_bram_77_tready),
        .ap_bram_77_addr0(ap_bram_iarg_77_addr0),
        .ap_bram_77_din0(ap_bram_iarg_77_din0),
        .ap_bram_77_dout0(ap_bram_iarg_77_dout0),
        .ap_bram_77_we0(ap_bram_iarg_77_we0),
        .ap_bram_77_en0(ap_bram_iarg_77_en0),
        .ap_bram_77_addr1(ap_bram_iarg_77_addr1),
        .ap_bram_77_din1(ap_bram_iarg_77_din1),
        .ap_bram_77_dout1(ap_bram_iarg_77_dout1),
        .ap_bram_77_we1(ap_bram_iarg_77_we1),
        .ap_bram_77_en1(ap_bram_iarg_77_en1),
        .s_axis_bram_78_tlast(s_axis_bram_78_tlast),
        .s_axis_bram_78_tvalid(s_axis_bram_78_tvalid),
        .s_axis_bram_78_tkeep(s_axis_bram_78_tkeep),
        .s_axis_bram_78_tstrb(s_axis_bram_78_tstrb),
        .s_axis_bram_78_tdata(s_axis_bram_78_tdata),
        .s_axis_bram_78_tready(s_axis_bram_78_tready),
        .ap_bram_78_addr0(ap_bram_iarg_78_addr0),
        .ap_bram_78_din0(ap_bram_iarg_78_din0),
        .ap_bram_78_dout0(ap_bram_iarg_78_dout0),
        .ap_bram_78_we0(ap_bram_iarg_78_we0),
        .ap_bram_78_en0(ap_bram_iarg_78_en0),
        .ap_bram_78_addr1(ap_bram_iarg_78_addr1),
        .ap_bram_78_din1(ap_bram_iarg_78_din1),
        .ap_bram_78_dout1(ap_bram_iarg_78_dout1),
        .ap_bram_78_we1(ap_bram_iarg_78_we1),
        .ap_bram_78_en1(ap_bram_iarg_78_en1),
        .s_axis_bram_79_tlast(s_axis_bram_79_tlast),
        .s_axis_bram_79_tvalid(s_axis_bram_79_tvalid),
        .s_axis_bram_79_tkeep(s_axis_bram_79_tkeep),
        .s_axis_bram_79_tstrb(s_axis_bram_79_tstrb),
        .s_axis_bram_79_tdata(s_axis_bram_79_tdata),
        .s_axis_bram_79_tready(s_axis_bram_79_tready),
        .ap_bram_79_addr0(ap_bram_iarg_79_addr0),
        .ap_bram_79_din0(ap_bram_iarg_79_din0),
        .ap_bram_79_dout0(ap_bram_iarg_79_dout0),
        .ap_bram_79_we0(ap_bram_iarg_79_we0),
        .ap_bram_79_en0(ap_bram_iarg_79_en0),
        .ap_bram_79_addr1(ap_bram_iarg_79_addr1),
        .ap_bram_79_din1(ap_bram_iarg_79_din1),
        .ap_bram_79_dout1(ap_bram_iarg_79_dout1),
        .ap_bram_79_we1(ap_bram_iarg_79_we1),
        .ap_bram_79_en1(ap_bram_iarg_79_en1),
        .s_axis_bram_80_tlast(s_axis_bram_80_tlast),
        .s_axis_bram_80_tvalid(s_axis_bram_80_tvalid),
        .s_axis_bram_80_tkeep(s_axis_bram_80_tkeep),
        .s_axis_bram_80_tstrb(s_axis_bram_80_tstrb),
        .s_axis_bram_80_tdata(s_axis_bram_80_tdata),
        .s_axis_bram_80_tready(s_axis_bram_80_tready),
        .ap_bram_80_addr0(ap_bram_iarg_80_addr0),
        .ap_bram_80_din0(ap_bram_iarg_80_din0),
        .ap_bram_80_dout0(ap_bram_iarg_80_dout0),
        .ap_bram_80_we0(ap_bram_iarg_80_we0),
        .ap_bram_80_en0(ap_bram_iarg_80_en0),
        .ap_bram_80_addr1(ap_bram_iarg_80_addr1),
        .ap_bram_80_din1(ap_bram_iarg_80_din1),
        .ap_bram_80_dout1(ap_bram_iarg_80_dout1),
        .ap_bram_80_we1(ap_bram_iarg_80_we1),
        .ap_bram_80_en1(ap_bram_iarg_80_en1),
        .s_axis_bram_81_tlast(s_axis_bram_81_tlast),
        .s_axis_bram_81_tvalid(s_axis_bram_81_tvalid),
        .s_axis_bram_81_tkeep(s_axis_bram_81_tkeep),
        .s_axis_bram_81_tstrb(s_axis_bram_81_tstrb),
        .s_axis_bram_81_tdata(s_axis_bram_81_tdata),
        .s_axis_bram_81_tready(s_axis_bram_81_tready),
        .ap_bram_81_addr0(ap_bram_iarg_81_addr0),
        .ap_bram_81_din0(ap_bram_iarg_81_din0),
        .ap_bram_81_dout0(ap_bram_iarg_81_dout0),
        .ap_bram_81_we0(ap_bram_iarg_81_we0),
        .ap_bram_81_en0(ap_bram_iarg_81_en0),
        .ap_bram_81_addr1(ap_bram_iarg_81_addr1),
        .ap_bram_81_din1(ap_bram_iarg_81_din1),
        .ap_bram_81_dout1(ap_bram_iarg_81_dout1),
        .ap_bram_81_we1(ap_bram_iarg_81_we1),
        .ap_bram_81_en1(ap_bram_iarg_81_en1),
        .s_axis_bram_82_tlast(s_axis_bram_82_tlast),
        .s_axis_bram_82_tvalid(s_axis_bram_82_tvalid),
        .s_axis_bram_82_tkeep(s_axis_bram_82_tkeep),
        .s_axis_bram_82_tstrb(s_axis_bram_82_tstrb),
        .s_axis_bram_82_tdata(s_axis_bram_82_tdata),
        .s_axis_bram_82_tready(s_axis_bram_82_tready),
        .ap_bram_82_addr0(ap_bram_iarg_82_addr0),
        .ap_bram_82_din0(ap_bram_iarg_82_din0),
        .ap_bram_82_dout0(ap_bram_iarg_82_dout0),
        .ap_bram_82_we0(ap_bram_iarg_82_we0),
        .ap_bram_82_en0(ap_bram_iarg_82_en0),
        .ap_bram_82_addr1(ap_bram_iarg_82_addr1),
        .ap_bram_82_din1(ap_bram_iarg_82_din1),
        .ap_bram_82_dout1(ap_bram_iarg_82_dout1),
        .ap_bram_82_we1(ap_bram_iarg_82_we1),
        .ap_bram_82_en1(ap_bram_iarg_82_en1),
        .s_axis_bram_83_tlast(s_axis_bram_83_tlast),
        .s_axis_bram_83_tvalid(s_axis_bram_83_tvalid),
        .s_axis_bram_83_tkeep(s_axis_bram_83_tkeep),
        .s_axis_bram_83_tstrb(s_axis_bram_83_tstrb),
        .s_axis_bram_83_tdata(s_axis_bram_83_tdata),
        .s_axis_bram_83_tready(s_axis_bram_83_tready),
        .ap_bram_83_addr0(ap_bram_iarg_83_addr0),
        .ap_bram_83_din0(ap_bram_iarg_83_din0),
        .ap_bram_83_dout0(ap_bram_iarg_83_dout0),
        .ap_bram_83_we0(ap_bram_iarg_83_we0),
        .ap_bram_83_en0(ap_bram_iarg_83_en0),
        .ap_bram_83_addr1(ap_bram_iarg_83_addr1),
        .ap_bram_83_din1(ap_bram_iarg_83_din1),
        .ap_bram_83_dout1(ap_bram_iarg_83_dout1),
        .ap_bram_83_we1(ap_bram_iarg_83_we1),
        .ap_bram_83_en1(ap_bram_iarg_83_en1),
        .s_axis_bram_84_tlast(s_axis_bram_84_tlast),
        .s_axis_bram_84_tvalid(s_axis_bram_84_tvalid),
        .s_axis_bram_84_tkeep(s_axis_bram_84_tkeep),
        .s_axis_bram_84_tstrb(s_axis_bram_84_tstrb),
        .s_axis_bram_84_tdata(s_axis_bram_84_tdata),
        .s_axis_bram_84_tready(s_axis_bram_84_tready),
        .ap_bram_84_addr0(ap_bram_iarg_84_addr0),
        .ap_bram_84_din0(ap_bram_iarg_84_din0),
        .ap_bram_84_dout0(ap_bram_iarg_84_dout0),
        .ap_bram_84_we0(ap_bram_iarg_84_we0),
        .ap_bram_84_en0(ap_bram_iarg_84_en0),
        .ap_bram_84_addr1(ap_bram_iarg_84_addr1),
        .ap_bram_84_din1(ap_bram_iarg_84_din1),
        .ap_bram_84_dout1(ap_bram_iarg_84_dout1),
        .ap_bram_84_we1(ap_bram_iarg_84_we1),
        .ap_bram_84_en1(ap_bram_iarg_84_en1),
        .s_axis_bram_85_tlast(s_axis_bram_85_tlast),
        .s_axis_bram_85_tvalid(s_axis_bram_85_tvalid),
        .s_axis_bram_85_tkeep(s_axis_bram_85_tkeep),
        .s_axis_bram_85_tstrb(s_axis_bram_85_tstrb),
        .s_axis_bram_85_tdata(s_axis_bram_85_tdata),
        .s_axis_bram_85_tready(s_axis_bram_85_tready),
        .ap_bram_85_addr0(ap_bram_iarg_85_addr0),
        .ap_bram_85_din0(ap_bram_iarg_85_din0),
        .ap_bram_85_dout0(ap_bram_iarg_85_dout0),
        .ap_bram_85_we0(ap_bram_iarg_85_we0),
        .ap_bram_85_en0(ap_bram_iarg_85_en0),
        .ap_bram_85_addr1(ap_bram_iarg_85_addr1),
        .ap_bram_85_din1(ap_bram_iarg_85_din1),
        .ap_bram_85_dout1(ap_bram_iarg_85_dout1),
        .ap_bram_85_we1(ap_bram_iarg_85_we1),
        .ap_bram_85_en1(ap_bram_iarg_85_en1),
        .s_axis_bram_86_tlast(s_axis_bram_86_tlast),
        .s_axis_bram_86_tvalid(s_axis_bram_86_tvalid),
        .s_axis_bram_86_tkeep(s_axis_bram_86_tkeep),
        .s_axis_bram_86_tstrb(s_axis_bram_86_tstrb),
        .s_axis_bram_86_tdata(s_axis_bram_86_tdata),
        .s_axis_bram_86_tready(s_axis_bram_86_tready),
        .ap_bram_86_addr0(ap_bram_iarg_86_addr0),
        .ap_bram_86_din0(ap_bram_iarg_86_din0),
        .ap_bram_86_dout0(ap_bram_iarg_86_dout0),
        .ap_bram_86_we0(ap_bram_iarg_86_we0),
        .ap_bram_86_en0(ap_bram_iarg_86_en0),
        .ap_bram_86_addr1(ap_bram_iarg_86_addr1),
        .ap_bram_86_din1(ap_bram_iarg_86_din1),
        .ap_bram_86_dout1(ap_bram_iarg_86_dout1),
        .ap_bram_86_we1(ap_bram_iarg_86_we1),
        .ap_bram_86_en1(ap_bram_iarg_86_en1),
        .s_axis_bram_87_tlast(s_axis_bram_87_tlast),
        .s_axis_bram_87_tvalid(s_axis_bram_87_tvalid),
        .s_axis_bram_87_tkeep(s_axis_bram_87_tkeep),
        .s_axis_bram_87_tstrb(s_axis_bram_87_tstrb),
        .s_axis_bram_87_tdata(s_axis_bram_87_tdata),
        .s_axis_bram_87_tready(s_axis_bram_87_tready),
        .ap_bram_87_addr0(ap_bram_iarg_87_addr0),
        .ap_bram_87_din0(ap_bram_iarg_87_din0),
        .ap_bram_87_dout0(ap_bram_iarg_87_dout0),
        .ap_bram_87_we0(ap_bram_iarg_87_we0),
        .ap_bram_87_en0(ap_bram_iarg_87_en0),
        .ap_bram_87_addr1(ap_bram_iarg_87_addr1),
        .ap_bram_87_din1(ap_bram_iarg_87_din1),
        .ap_bram_87_dout1(ap_bram_iarg_87_dout1),
        .ap_bram_87_we1(ap_bram_iarg_87_we1),
        .ap_bram_87_en1(ap_bram_iarg_87_en1),
        .s_axis_bram_88_tlast(s_axis_bram_88_tlast),
        .s_axis_bram_88_tvalid(s_axis_bram_88_tvalid),
        .s_axis_bram_88_tkeep(s_axis_bram_88_tkeep),
        .s_axis_bram_88_tstrb(s_axis_bram_88_tstrb),
        .s_axis_bram_88_tdata(s_axis_bram_88_tdata),
        .s_axis_bram_88_tready(s_axis_bram_88_tready),
        .ap_bram_88_addr0(ap_bram_iarg_88_addr0),
        .ap_bram_88_din0(ap_bram_iarg_88_din0),
        .ap_bram_88_dout0(ap_bram_iarg_88_dout0),
        .ap_bram_88_we0(ap_bram_iarg_88_we0),
        .ap_bram_88_en0(ap_bram_iarg_88_en0),
        .ap_bram_88_addr1(ap_bram_iarg_88_addr1),
        .ap_bram_88_din1(ap_bram_iarg_88_din1),
        .ap_bram_88_dout1(ap_bram_iarg_88_dout1),
        .ap_bram_88_we1(ap_bram_iarg_88_we1),
        .ap_bram_88_en1(ap_bram_iarg_88_en1),
        .s_axis_bram_89_tlast(s_axis_bram_89_tlast),
        .s_axis_bram_89_tvalid(s_axis_bram_89_tvalid),
        .s_axis_bram_89_tkeep(s_axis_bram_89_tkeep),
        .s_axis_bram_89_tstrb(s_axis_bram_89_tstrb),
        .s_axis_bram_89_tdata(s_axis_bram_89_tdata),
        .s_axis_bram_89_tready(s_axis_bram_89_tready),
        .ap_bram_89_addr0(ap_bram_iarg_89_addr0),
        .ap_bram_89_din0(ap_bram_iarg_89_din0),
        .ap_bram_89_dout0(ap_bram_iarg_89_dout0),
        .ap_bram_89_we0(ap_bram_iarg_89_we0),
        .ap_bram_89_en0(ap_bram_iarg_89_en0),
        .ap_bram_89_addr1(ap_bram_iarg_89_addr1),
        .ap_bram_89_din1(ap_bram_iarg_89_din1),
        .ap_bram_89_dout1(ap_bram_iarg_89_dout1),
        .ap_bram_89_we1(ap_bram_iarg_89_we1),
        .ap_bram_89_en1(ap_bram_iarg_89_en1),
        .s_axis_bram_90_tlast(s_axis_bram_90_tlast),
        .s_axis_bram_90_tvalid(s_axis_bram_90_tvalid),
        .s_axis_bram_90_tkeep(s_axis_bram_90_tkeep),
        .s_axis_bram_90_tstrb(s_axis_bram_90_tstrb),
        .s_axis_bram_90_tdata(s_axis_bram_90_tdata),
        .s_axis_bram_90_tready(s_axis_bram_90_tready),
        .ap_bram_90_addr0(ap_bram_iarg_90_addr0),
        .ap_bram_90_din0(ap_bram_iarg_90_din0),
        .ap_bram_90_dout0(ap_bram_iarg_90_dout0),
        .ap_bram_90_we0(ap_bram_iarg_90_we0),
        .ap_bram_90_en0(ap_bram_iarg_90_en0),
        .ap_bram_90_addr1(ap_bram_iarg_90_addr1),
        .ap_bram_90_din1(ap_bram_iarg_90_din1),
        .ap_bram_90_dout1(ap_bram_iarg_90_dout1),
        .ap_bram_90_we1(ap_bram_iarg_90_we1),
        .ap_bram_90_en1(ap_bram_iarg_90_en1),
        .s_axis_bram_91_tlast(s_axis_bram_91_tlast),
        .s_axis_bram_91_tvalid(s_axis_bram_91_tvalid),
        .s_axis_bram_91_tkeep(s_axis_bram_91_tkeep),
        .s_axis_bram_91_tstrb(s_axis_bram_91_tstrb),
        .s_axis_bram_91_tdata(s_axis_bram_91_tdata),
        .s_axis_bram_91_tready(s_axis_bram_91_tready),
        .ap_bram_91_addr0(ap_bram_iarg_91_addr0),
        .ap_bram_91_din0(ap_bram_iarg_91_din0),
        .ap_bram_91_dout0(ap_bram_iarg_91_dout0),
        .ap_bram_91_we0(ap_bram_iarg_91_we0),
        .ap_bram_91_en0(ap_bram_iarg_91_en0),
        .ap_bram_91_addr1(ap_bram_iarg_91_addr1),
        .ap_bram_91_din1(ap_bram_iarg_91_din1),
        .ap_bram_91_dout1(ap_bram_iarg_91_dout1),
        .ap_bram_91_we1(ap_bram_iarg_91_we1),
        .ap_bram_91_en1(ap_bram_iarg_91_en1),
        .s_axis_bram_92_tlast(s_axis_bram_92_tlast),
        .s_axis_bram_92_tvalid(s_axis_bram_92_tvalid),
        .s_axis_bram_92_tkeep(s_axis_bram_92_tkeep),
        .s_axis_bram_92_tstrb(s_axis_bram_92_tstrb),
        .s_axis_bram_92_tdata(s_axis_bram_92_tdata),
        .s_axis_bram_92_tready(s_axis_bram_92_tready),
        .ap_bram_92_addr0(ap_bram_iarg_92_addr0),
        .ap_bram_92_din0(ap_bram_iarg_92_din0),
        .ap_bram_92_dout0(ap_bram_iarg_92_dout0),
        .ap_bram_92_we0(ap_bram_iarg_92_we0),
        .ap_bram_92_en0(ap_bram_iarg_92_en0),
        .ap_bram_92_addr1(ap_bram_iarg_92_addr1),
        .ap_bram_92_din1(ap_bram_iarg_92_din1),
        .ap_bram_92_dout1(ap_bram_iarg_92_dout1),
        .ap_bram_92_we1(ap_bram_iarg_92_we1),
        .ap_bram_92_en1(ap_bram_iarg_92_en1),
        .s_axis_bram_93_tlast(s_axis_bram_93_tlast),
        .s_axis_bram_93_tvalid(s_axis_bram_93_tvalid),
        .s_axis_bram_93_tkeep(s_axis_bram_93_tkeep),
        .s_axis_bram_93_tstrb(s_axis_bram_93_tstrb),
        .s_axis_bram_93_tdata(s_axis_bram_93_tdata),
        .s_axis_bram_93_tready(s_axis_bram_93_tready),
        .ap_bram_93_addr0(ap_bram_iarg_93_addr0),
        .ap_bram_93_din0(ap_bram_iarg_93_din0),
        .ap_bram_93_dout0(ap_bram_iarg_93_dout0),
        .ap_bram_93_we0(ap_bram_iarg_93_we0),
        .ap_bram_93_en0(ap_bram_iarg_93_en0),
        .ap_bram_93_addr1(ap_bram_iarg_93_addr1),
        .ap_bram_93_din1(ap_bram_iarg_93_din1),
        .ap_bram_93_dout1(ap_bram_iarg_93_dout1),
        .ap_bram_93_we1(ap_bram_iarg_93_we1),
        .ap_bram_93_en1(ap_bram_iarg_93_en1),
        .s_axis_bram_94_tlast(s_axis_bram_94_tlast),
        .s_axis_bram_94_tvalid(s_axis_bram_94_tvalid),
        .s_axis_bram_94_tkeep(s_axis_bram_94_tkeep),
        .s_axis_bram_94_tstrb(s_axis_bram_94_tstrb),
        .s_axis_bram_94_tdata(s_axis_bram_94_tdata),
        .s_axis_bram_94_tready(s_axis_bram_94_tready),
        .ap_bram_94_addr0(ap_bram_iarg_94_addr0),
        .ap_bram_94_din0(ap_bram_iarg_94_din0),
        .ap_bram_94_dout0(ap_bram_iarg_94_dout0),
        .ap_bram_94_we0(ap_bram_iarg_94_we0),
        .ap_bram_94_en0(ap_bram_iarg_94_en0),
        .ap_bram_94_addr1(ap_bram_iarg_94_addr1),
        .ap_bram_94_din1(ap_bram_iarg_94_din1),
        .ap_bram_94_dout1(ap_bram_iarg_94_dout1),
        .ap_bram_94_we1(ap_bram_iarg_94_we1),
        .ap_bram_94_en1(ap_bram_iarg_94_en1),
        .s_axis_bram_95_tlast(s_axis_bram_95_tlast),
        .s_axis_bram_95_tvalid(s_axis_bram_95_tvalid),
        .s_axis_bram_95_tkeep(s_axis_bram_95_tkeep),
        .s_axis_bram_95_tstrb(s_axis_bram_95_tstrb),
        .s_axis_bram_95_tdata(s_axis_bram_95_tdata),
        .s_axis_bram_95_tready(s_axis_bram_95_tready),
        .ap_bram_95_addr0(ap_bram_iarg_95_addr0),
        .ap_bram_95_din0(ap_bram_iarg_95_din0),
        .ap_bram_95_dout0(ap_bram_iarg_95_dout0),
        .ap_bram_95_we0(ap_bram_iarg_95_we0),
        .ap_bram_95_en0(ap_bram_iarg_95_en0),
        .ap_bram_95_addr1(ap_bram_iarg_95_addr1),
        .ap_bram_95_din1(ap_bram_iarg_95_din1),
        .ap_bram_95_dout1(ap_bram_iarg_95_dout1),
        .ap_bram_95_we1(ap_bram_iarg_95_we1),
        .ap_bram_95_en1(ap_bram_iarg_95_en1),
        .s_axis_bram_96_tlast(s_axis_bram_96_tlast),
        .s_axis_bram_96_tvalid(s_axis_bram_96_tvalid),
        .s_axis_bram_96_tkeep(s_axis_bram_96_tkeep),
        .s_axis_bram_96_tstrb(s_axis_bram_96_tstrb),
        .s_axis_bram_96_tdata(s_axis_bram_96_tdata),
        .s_axis_bram_96_tready(s_axis_bram_96_tready),
        .ap_bram_96_addr0(ap_bram_iarg_96_addr0),
        .ap_bram_96_din0(ap_bram_iarg_96_din0),
        .ap_bram_96_dout0(ap_bram_iarg_96_dout0),
        .ap_bram_96_we0(ap_bram_iarg_96_we0),
        .ap_bram_96_en0(ap_bram_iarg_96_en0),
        .ap_bram_96_addr1(ap_bram_iarg_96_addr1),
        .ap_bram_96_din1(ap_bram_iarg_96_din1),
        .ap_bram_96_dout1(ap_bram_iarg_96_dout1),
        .ap_bram_96_we1(ap_bram_iarg_96_we1),
        .ap_bram_96_en1(ap_bram_iarg_96_en1),
        .s_axis_bram_97_tlast(s_axis_bram_97_tlast),
        .s_axis_bram_97_tvalid(s_axis_bram_97_tvalid),
        .s_axis_bram_97_tkeep(s_axis_bram_97_tkeep),
        .s_axis_bram_97_tstrb(s_axis_bram_97_tstrb),
        .s_axis_bram_97_tdata(s_axis_bram_97_tdata),
        .s_axis_bram_97_tready(s_axis_bram_97_tready),
        .ap_bram_97_addr0(ap_bram_iarg_97_addr0),
        .ap_bram_97_din0(ap_bram_iarg_97_din0),
        .ap_bram_97_dout0(ap_bram_iarg_97_dout0),
        .ap_bram_97_we0(ap_bram_iarg_97_we0),
        .ap_bram_97_en0(ap_bram_iarg_97_en0),
        .ap_bram_97_addr1(ap_bram_iarg_97_addr1),
        .ap_bram_97_din1(ap_bram_iarg_97_din1),
        .ap_bram_97_dout1(ap_bram_iarg_97_dout1),
        .ap_bram_97_we1(ap_bram_iarg_97_we1),
        .ap_bram_97_en1(ap_bram_iarg_97_en1),
        .s_axis_bram_98_tlast(s_axis_bram_98_tlast),
        .s_axis_bram_98_tvalid(s_axis_bram_98_tvalid),
        .s_axis_bram_98_tkeep(s_axis_bram_98_tkeep),
        .s_axis_bram_98_tstrb(s_axis_bram_98_tstrb),
        .s_axis_bram_98_tdata(s_axis_bram_98_tdata),
        .s_axis_bram_98_tready(s_axis_bram_98_tready),
        .ap_bram_98_addr0(ap_bram_iarg_98_addr0),
        .ap_bram_98_din0(ap_bram_iarg_98_din0),
        .ap_bram_98_dout0(ap_bram_iarg_98_dout0),
        .ap_bram_98_we0(ap_bram_iarg_98_we0),
        .ap_bram_98_en0(ap_bram_iarg_98_en0),
        .ap_bram_98_addr1(ap_bram_iarg_98_addr1),
        .ap_bram_98_din1(ap_bram_iarg_98_din1),
        .ap_bram_98_dout1(ap_bram_iarg_98_dout1),
        .ap_bram_98_we1(ap_bram_iarg_98_we1),
        .ap_bram_98_en1(ap_bram_iarg_98_en1),
        .s_axis_bram_99_tlast(s_axis_bram_99_tlast),
        .s_axis_bram_99_tvalid(s_axis_bram_99_tvalid),
        .s_axis_bram_99_tkeep(s_axis_bram_99_tkeep),
        .s_axis_bram_99_tstrb(s_axis_bram_99_tstrb),
        .s_axis_bram_99_tdata(s_axis_bram_99_tdata),
        .s_axis_bram_99_tready(s_axis_bram_99_tready),
        .ap_bram_99_addr0(ap_bram_iarg_99_addr0),
        .ap_bram_99_din0(ap_bram_iarg_99_din0),
        .ap_bram_99_dout0(ap_bram_iarg_99_dout0),
        .ap_bram_99_we0(ap_bram_iarg_99_we0),
        .ap_bram_99_en0(ap_bram_iarg_99_en0),
        .ap_bram_99_addr1(ap_bram_iarg_99_addr1),
        .ap_bram_99_din1(ap_bram_iarg_99_din1),
        .ap_bram_99_dout1(ap_bram_iarg_99_dout1),
        .ap_bram_99_we1(ap_bram_iarg_99_we1),
        .ap_bram_99_en1(ap_bram_iarg_99_en1),
        .s_axis_bram_100_tlast(s_axis_bram_100_tlast),
        .s_axis_bram_100_tvalid(s_axis_bram_100_tvalid),
        .s_axis_bram_100_tkeep(s_axis_bram_100_tkeep),
        .s_axis_bram_100_tstrb(s_axis_bram_100_tstrb),
        .s_axis_bram_100_tdata(s_axis_bram_100_tdata),
        .s_axis_bram_100_tready(s_axis_bram_100_tready),
        .ap_bram_100_addr0(ap_bram_iarg_100_addr0),
        .ap_bram_100_din0(ap_bram_iarg_100_din0),
        .ap_bram_100_dout0(ap_bram_iarg_100_dout0),
        .ap_bram_100_we0(ap_bram_iarg_100_we0),
        .ap_bram_100_en0(ap_bram_iarg_100_en0),
        .ap_bram_100_addr1(ap_bram_iarg_100_addr1),
        .ap_bram_100_din1(ap_bram_iarg_100_din1),
        .ap_bram_100_dout1(ap_bram_iarg_100_dout1),
        .ap_bram_100_we1(ap_bram_iarg_100_we1),
        .ap_bram_100_en1(ap_bram_iarg_100_en1),
        .s_axis_bram_101_tlast(s_axis_bram_101_tlast),
        .s_axis_bram_101_tvalid(s_axis_bram_101_tvalid),
        .s_axis_bram_101_tkeep(s_axis_bram_101_tkeep),
        .s_axis_bram_101_tstrb(s_axis_bram_101_tstrb),
        .s_axis_bram_101_tdata(s_axis_bram_101_tdata),
        .s_axis_bram_101_tready(s_axis_bram_101_tready),
        .ap_bram_101_addr0(ap_bram_iarg_101_addr0),
        .ap_bram_101_din0(ap_bram_iarg_101_din0),
        .ap_bram_101_dout0(ap_bram_iarg_101_dout0),
        .ap_bram_101_we0(ap_bram_iarg_101_we0),
        .ap_bram_101_en0(ap_bram_iarg_101_en0),
        .ap_bram_101_addr1(ap_bram_iarg_101_addr1),
        .ap_bram_101_din1(ap_bram_iarg_101_din1),
        .ap_bram_101_dout1(ap_bram_iarg_101_dout1),
        .ap_bram_101_we1(ap_bram_iarg_101_we1),
        .ap_bram_101_en1(ap_bram_iarg_101_en1),
        .s_axis_bram_102_tlast(s_axis_bram_102_tlast),
        .s_axis_bram_102_tvalid(s_axis_bram_102_tvalid),
        .s_axis_bram_102_tkeep(s_axis_bram_102_tkeep),
        .s_axis_bram_102_tstrb(s_axis_bram_102_tstrb),
        .s_axis_bram_102_tdata(s_axis_bram_102_tdata),
        .s_axis_bram_102_tready(s_axis_bram_102_tready),
        .ap_bram_102_addr0(ap_bram_iarg_102_addr0),
        .ap_bram_102_din0(ap_bram_iarg_102_din0),
        .ap_bram_102_dout0(ap_bram_iarg_102_dout0),
        .ap_bram_102_we0(ap_bram_iarg_102_we0),
        .ap_bram_102_en0(ap_bram_iarg_102_en0),
        .ap_bram_102_addr1(ap_bram_iarg_102_addr1),
        .ap_bram_102_din1(ap_bram_iarg_102_din1),
        .ap_bram_102_dout1(ap_bram_iarg_102_dout1),
        .ap_bram_102_we1(ap_bram_iarg_102_we1),
        .ap_bram_102_en1(ap_bram_iarg_102_en1),
        .s_axis_bram_103_tlast(s_axis_bram_103_tlast),
        .s_axis_bram_103_tvalid(s_axis_bram_103_tvalid),
        .s_axis_bram_103_tkeep(s_axis_bram_103_tkeep),
        .s_axis_bram_103_tstrb(s_axis_bram_103_tstrb),
        .s_axis_bram_103_tdata(s_axis_bram_103_tdata),
        .s_axis_bram_103_tready(s_axis_bram_103_tready),
        .ap_bram_103_addr0(ap_bram_iarg_103_addr0),
        .ap_bram_103_din0(ap_bram_iarg_103_din0),
        .ap_bram_103_dout0(ap_bram_iarg_103_dout0),
        .ap_bram_103_we0(ap_bram_iarg_103_we0),
        .ap_bram_103_en0(ap_bram_iarg_103_en0),
        .ap_bram_103_addr1(ap_bram_iarg_103_addr1),
        .ap_bram_103_din1(ap_bram_iarg_103_din1),
        .ap_bram_103_dout1(ap_bram_iarg_103_dout1),
        .ap_bram_103_we1(ap_bram_iarg_103_we1),
        .ap_bram_103_en1(ap_bram_iarg_103_en1),
        .s_axis_bram_104_tlast(s_axis_bram_104_tlast),
        .s_axis_bram_104_tvalid(s_axis_bram_104_tvalid),
        .s_axis_bram_104_tkeep(s_axis_bram_104_tkeep),
        .s_axis_bram_104_tstrb(s_axis_bram_104_tstrb),
        .s_axis_bram_104_tdata(s_axis_bram_104_tdata),
        .s_axis_bram_104_tready(s_axis_bram_104_tready),
        .ap_bram_104_addr0(ap_bram_iarg_104_addr0),
        .ap_bram_104_din0(ap_bram_iarg_104_din0),
        .ap_bram_104_dout0(ap_bram_iarg_104_dout0),
        .ap_bram_104_we0(ap_bram_iarg_104_we0),
        .ap_bram_104_en0(ap_bram_iarg_104_en0),
        .ap_bram_104_addr1(ap_bram_iarg_104_addr1),
        .ap_bram_104_din1(ap_bram_iarg_104_din1),
        .ap_bram_104_dout1(ap_bram_iarg_104_dout1),
        .ap_bram_104_we1(ap_bram_iarg_104_we1),
        .ap_bram_104_en1(ap_bram_iarg_104_en1),
        .s_axis_bram_105_tlast(s_axis_bram_105_tlast),
        .s_axis_bram_105_tvalid(s_axis_bram_105_tvalid),
        .s_axis_bram_105_tkeep(s_axis_bram_105_tkeep),
        .s_axis_bram_105_tstrb(s_axis_bram_105_tstrb),
        .s_axis_bram_105_tdata(s_axis_bram_105_tdata),
        .s_axis_bram_105_tready(s_axis_bram_105_tready),
        .ap_bram_105_addr0(ap_bram_iarg_105_addr0),
        .ap_bram_105_din0(ap_bram_iarg_105_din0),
        .ap_bram_105_dout0(ap_bram_iarg_105_dout0),
        .ap_bram_105_we0(ap_bram_iarg_105_we0),
        .ap_bram_105_en0(ap_bram_iarg_105_en0),
        .ap_bram_105_addr1(ap_bram_iarg_105_addr1),
        .ap_bram_105_din1(ap_bram_iarg_105_din1),
        .ap_bram_105_dout1(ap_bram_iarg_105_dout1),
        .ap_bram_105_we1(ap_bram_iarg_105_we1),
        .ap_bram_105_en1(ap_bram_iarg_105_en1),
        .s_axis_bram_106_tlast(s_axis_bram_106_tlast),
        .s_axis_bram_106_tvalid(s_axis_bram_106_tvalid),
        .s_axis_bram_106_tkeep(s_axis_bram_106_tkeep),
        .s_axis_bram_106_tstrb(s_axis_bram_106_tstrb),
        .s_axis_bram_106_tdata(s_axis_bram_106_tdata),
        .s_axis_bram_106_tready(s_axis_bram_106_tready),
        .ap_bram_106_addr0(ap_bram_iarg_106_addr0),
        .ap_bram_106_din0(ap_bram_iarg_106_din0),
        .ap_bram_106_dout0(ap_bram_iarg_106_dout0),
        .ap_bram_106_we0(ap_bram_iarg_106_we0),
        .ap_bram_106_en0(ap_bram_iarg_106_en0),
        .ap_bram_106_addr1(ap_bram_iarg_106_addr1),
        .ap_bram_106_din1(ap_bram_iarg_106_din1),
        .ap_bram_106_dout1(ap_bram_iarg_106_dout1),
        .ap_bram_106_we1(ap_bram_iarg_106_we1),
        .ap_bram_106_en1(ap_bram_iarg_106_en1),
        .s_axis_bram_107_tlast(s_axis_bram_107_tlast),
        .s_axis_bram_107_tvalid(s_axis_bram_107_tvalid),
        .s_axis_bram_107_tkeep(s_axis_bram_107_tkeep),
        .s_axis_bram_107_tstrb(s_axis_bram_107_tstrb),
        .s_axis_bram_107_tdata(s_axis_bram_107_tdata),
        .s_axis_bram_107_tready(s_axis_bram_107_tready),
        .ap_bram_107_addr0(ap_bram_iarg_107_addr0),
        .ap_bram_107_din0(ap_bram_iarg_107_din0),
        .ap_bram_107_dout0(ap_bram_iarg_107_dout0),
        .ap_bram_107_we0(ap_bram_iarg_107_we0),
        .ap_bram_107_en0(ap_bram_iarg_107_en0),
        .ap_bram_107_addr1(ap_bram_iarg_107_addr1),
        .ap_bram_107_din1(ap_bram_iarg_107_din1),
        .ap_bram_107_dout1(ap_bram_iarg_107_dout1),
        .ap_bram_107_we1(ap_bram_iarg_107_we1),
        .ap_bram_107_en1(ap_bram_iarg_107_en1),
        .s_axis_bram_108_tlast(s_axis_bram_108_tlast),
        .s_axis_bram_108_tvalid(s_axis_bram_108_tvalid),
        .s_axis_bram_108_tkeep(s_axis_bram_108_tkeep),
        .s_axis_bram_108_tstrb(s_axis_bram_108_tstrb),
        .s_axis_bram_108_tdata(s_axis_bram_108_tdata),
        .s_axis_bram_108_tready(s_axis_bram_108_tready),
        .ap_bram_108_addr0(ap_bram_iarg_108_addr0),
        .ap_bram_108_din0(ap_bram_iarg_108_din0),
        .ap_bram_108_dout0(ap_bram_iarg_108_dout0),
        .ap_bram_108_we0(ap_bram_iarg_108_we0),
        .ap_bram_108_en0(ap_bram_iarg_108_en0),
        .ap_bram_108_addr1(ap_bram_iarg_108_addr1),
        .ap_bram_108_din1(ap_bram_iarg_108_din1),
        .ap_bram_108_dout1(ap_bram_iarg_108_dout1),
        .ap_bram_108_we1(ap_bram_iarg_108_we1),
        .ap_bram_108_en1(ap_bram_iarg_108_en1),
        .s_axis_bram_109_tlast(s_axis_bram_109_tlast),
        .s_axis_bram_109_tvalid(s_axis_bram_109_tvalid),
        .s_axis_bram_109_tkeep(s_axis_bram_109_tkeep),
        .s_axis_bram_109_tstrb(s_axis_bram_109_tstrb),
        .s_axis_bram_109_tdata(s_axis_bram_109_tdata),
        .s_axis_bram_109_tready(s_axis_bram_109_tready),
        .ap_bram_109_addr0(ap_bram_iarg_109_addr0),
        .ap_bram_109_din0(ap_bram_iarg_109_din0),
        .ap_bram_109_dout0(ap_bram_iarg_109_dout0),
        .ap_bram_109_we0(ap_bram_iarg_109_we0),
        .ap_bram_109_en0(ap_bram_iarg_109_en0),
        .ap_bram_109_addr1(ap_bram_iarg_109_addr1),
        .ap_bram_109_din1(ap_bram_iarg_109_din1),
        .ap_bram_109_dout1(ap_bram_iarg_109_dout1),
        .ap_bram_109_we1(ap_bram_iarg_109_we1),
        .ap_bram_109_en1(ap_bram_iarg_109_en1),
        .s_axis_bram_110_tlast(s_axis_bram_110_tlast),
        .s_axis_bram_110_tvalid(s_axis_bram_110_tvalid),
        .s_axis_bram_110_tkeep(s_axis_bram_110_tkeep),
        .s_axis_bram_110_tstrb(s_axis_bram_110_tstrb),
        .s_axis_bram_110_tdata(s_axis_bram_110_tdata),
        .s_axis_bram_110_tready(s_axis_bram_110_tready),
        .ap_bram_110_addr0(ap_bram_iarg_110_addr0),
        .ap_bram_110_din0(ap_bram_iarg_110_din0),
        .ap_bram_110_dout0(ap_bram_iarg_110_dout0),
        .ap_bram_110_we0(ap_bram_iarg_110_we0),
        .ap_bram_110_en0(ap_bram_iarg_110_en0),
        .ap_bram_110_addr1(ap_bram_iarg_110_addr1),
        .ap_bram_110_din1(ap_bram_iarg_110_din1),
        .ap_bram_110_dout1(ap_bram_iarg_110_dout1),
        .ap_bram_110_we1(ap_bram_iarg_110_we1),
        .ap_bram_110_en1(ap_bram_iarg_110_en1),
        .s_axis_bram_111_tlast(s_axis_bram_111_tlast),
        .s_axis_bram_111_tvalid(s_axis_bram_111_tvalid),
        .s_axis_bram_111_tkeep(s_axis_bram_111_tkeep),
        .s_axis_bram_111_tstrb(s_axis_bram_111_tstrb),
        .s_axis_bram_111_tdata(s_axis_bram_111_tdata),
        .s_axis_bram_111_tready(s_axis_bram_111_tready),
        .ap_bram_111_addr0(ap_bram_iarg_111_addr0),
        .ap_bram_111_din0(ap_bram_iarg_111_din0),
        .ap_bram_111_dout0(ap_bram_iarg_111_dout0),
        .ap_bram_111_we0(ap_bram_iarg_111_we0),
        .ap_bram_111_en0(ap_bram_iarg_111_en0),
        .ap_bram_111_addr1(ap_bram_iarg_111_addr1),
        .ap_bram_111_din1(ap_bram_iarg_111_din1),
        .ap_bram_111_dout1(ap_bram_iarg_111_dout1),
        .ap_bram_111_we1(ap_bram_iarg_111_we1),
        .ap_bram_111_en1(ap_bram_iarg_111_en1),
        .s_axis_bram_112_tlast(s_axis_bram_112_tlast),
        .s_axis_bram_112_tvalid(s_axis_bram_112_tvalid),
        .s_axis_bram_112_tkeep(s_axis_bram_112_tkeep),
        .s_axis_bram_112_tstrb(s_axis_bram_112_tstrb),
        .s_axis_bram_112_tdata(s_axis_bram_112_tdata),
        .s_axis_bram_112_tready(s_axis_bram_112_tready),
        .ap_bram_112_addr0(ap_bram_iarg_112_addr0),
        .ap_bram_112_din0(ap_bram_iarg_112_din0),
        .ap_bram_112_dout0(ap_bram_iarg_112_dout0),
        .ap_bram_112_we0(ap_bram_iarg_112_we0),
        .ap_bram_112_en0(ap_bram_iarg_112_en0),
        .ap_bram_112_addr1(ap_bram_iarg_112_addr1),
        .ap_bram_112_din1(ap_bram_iarg_112_din1),
        .ap_bram_112_dout1(ap_bram_iarg_112_dout1),
        .ap_bram_112_we1(ap_bram_iarg_112_we1),
        .ap_bram_112_en1(ap_bram_iarg_112_en1),
        .s_axis_bram_113_tlast(s_axis_bram_113_tlast),
        .s_axis_bram_113_tvalid(s_axis_bram_113_tvalid),
        .s_axis_bram_113_tkeep(s_axis_bram_113_tkeep),
        .s_axis_bram_113_tstrb(s_axis_bram_113_tstrb),
        .s_axis_bram_113_tdata(s_axis_bram_113_tdata),
        .s_axis_bram_113_tready(s_axis_bram_113_tready),
        .ap_bram_113_addr0(ap_bram_iarg_113_addr0),
        .ap_bram_113_din0(ap_bram_iarg_113_din0),
        .ap_bram_113_dout0(ap_bram_iarg_113_dout0),
        .ap_bram_113_we0(ap_bram_iarg_113_we0),
        .ap_bram_113_en0(ap_bram_iarg_113_en0),
        .ap_bram_113_addr1(ap_bram_iarg_113_addr1),
        .ap_bram_113_din1(ap_bram_iarg_113_din1),
        .ap_bram_113_dout1(ap_bram_iarg_113_dout1),
        .ap_bram_113_we1(ap_bram_iarg_113_we1),
        .ap_bram_113_en1(ap_bram_iarg_113_en1),
        .s_axis_bram_114_tlast(s_axis_bram_114_tlast),
        .s_axis_bram_114_tvalid(s_axis_bram_114_tvalid),
        .s_axis_bram_114_tkeep(s_axis_bram_114_tkeep),
        .s_axis_bram_114_tstrb(s_axis_bram_114_tstrb),
        .s_axis_bram_114_tdata(s_axis_bram_114_tdata),
        .s_axis_bram_114_tready(s_axis_bram_114_tready),
        .ap_bram_114_addr0(ap_bram_iarg_114_addr0),
        .ap_bram_114_din0(ap_bram_iarg_114_din0),
        .ap_bram_114_dout0(ap_bram_iarg_114_dout0),
        .ap_bram_114_we0(ap_bram_iarg_114_we0),
        .ap_bram_114_en0(ap_bram_iarg_114_en0),
        .ap_bram_114_addr1(ap_bram_iarg_114_addr1),
        .ap_bram_114_din1(ap_bram_iarg_114_din1),
        .ap_bram_114_dout1(ap_bram_iarg_114_dout1),
        .ap_bram_114_we1(ap_bram_iarg_114_we1),
        .ap_bram_114_en1(ap_bram_iarg_114_en1),
        .s_axis_bram_115_tlast(s_axis_bram_115_tlast),
        .s_axis_bram_115_tvalid(s_axis_bram_115_tvalid),
        .s_axis_bram_115_tkeep(s_axis_bram_115_tkeep),
        .s_axis_bram_115_tstrb(s_axis_bram_115_tstrb),
        .s_axis_bram_115_tdata(s_axis_bram_115_tdata),
        .s_axis_bram_115_tready(s_axis_bram_115_tready),
        .ap_bram_115_addr0(ap_bram_iarg_115_addr0),
        .ap_bram_115_din0(ap_bram_iarg_115_din0),
        .ap_bram_115_dout0(ap_bram_iarg_115_dout0),
        .ap_bram_115_we0(ap_bram_iarg_115_we0),
        .ap_bram_115_en0(ap_bram_iarg_115_en0),
        .ap_bram_115_addr1(ap_bram_iarg_115_addr1),
        .ap_bram_115_din1(ap_bram_iarg_115_din1),
        .ap_bram_115_dout1(ap_bram_iarg_115_dout1),
        .ap_bram_115_we1(ap_bram_iarg_115_we1),
        .ap_bram_115_en1(ap_bram_iarg_115_en1),
        .s_axis_bram_116_tlast(s_axis_bram_116_tlast),
        .s_axis_bram_116_tvalid(s_axis_bram_116_tvalid),
        .s_axis_bram_116_tkeep(s_axis_bram_116_tkeep),
        .s_axis_bram_116_tstrb(s_axis_bram_116_tstrb),
        .s_axis_bram_116_tdata(s_axis_bram_116_tdata),
        .s_axis_bram_116_tready(s_axis_bram_116_tready),
        .ap_bram_116_addr0(ap_bram_iarg_116_addr0),
        .ap_bram_116_din0(ap_bram_iarg_116_din0),
        .ap_bram_116_dout0(ap_bram_iarg_116_dout0),
        .ap_bram_116_we0(ap_bram_iarg_116_we0),
        .ap_bram_116_en0(ap_bram_iarg_116_en0),
        .ap_bram_116_addr1(ap_bram_iarg_116_addr1),
        .ap_bram_116_din1(ap_bram_iarg_116_din1),
        .ap_bram_116_dout1(ap_bram_iarg_116_dout1),
        .ap_bram_116_we1(ap_bram_iarg_116_we1),
        .ap_bram_116_en1(ap_bram_iarg_116_en1),
        .s_axis_bram_117_tlast(s_axis_bram_117_tlast),
        .s_axis_bram_117_tvalid(s_axis_bram_117_tvalid),
        .s_axis_bram_117_tkeep(s_axis_bram_117_tkeep),
        .s_axis_bram_117_tstrb(s_axis_bram_117_tstrb),
        .s_axis_bram_117_tdata(s_axis_bram_117_tdata),
        .s_axis_bram_117_tready(s_axis_bram_117_tready),
        .ap_bram_117_addr0(ap_bram_iarg_117_addr0),
        .ap_bram_117_din0(ap_bram_iarg_117_din0),
        .ap_bram_117_dout0(ap_bram_iarg_117_dout0),
        .ap_bram_117_we0(ap_bram_iarg_117_we0),
        .ap_bram_117_en0(ap_bram_iarg_117_en0),
        .ap_bram_117_addr1(ap_bram_iarg_117_addr1),
        .ap_bram_117_din1(ap_bram_iarg_117_din1),
        .ap_bram_117_dout1(ap_bram_iarg_117_dout1),
        .ap_bram_117_we1(ap_bram_iarg_117_we1),
        .ap_bram_117_en1(ap_bram_iarg_117_en1),
        .s_axis_bram_118_tlast(s_axis_bram_118_tlast),
        .s_axis_bram_118_tvalid(s_axis_bram_118_tvalid),
        .s_axis_bram_118_tkeep(s_axis_bram_118_tkeep),
        .s_axis_bram_118_tstrb(s_axis_bram_118_tstrb),
        .s_axis_bram_118_tdata(s_axis_bram_118_tdata),
        .s_axis_bram_118_tready(s_axis_bram_118_tready),
        .ap_bram_118_addr0(ap_bram_iarg_118_addr0),
        .ap_bram_118_din0(ap_bram_iarg_118_din0),
        .ap_bram_118_dout0(ap_bram_iarg_118_dout0),
        .ap_bram_118_we0(ap_bram_iarg_118_we0),
        .ap_bram_118_en0(ap_bram_iarg_118_en0),
        .ap_bram_118_addr1(ap_bram_iarg_118_addr1),
        .ap_bram_118_din1(ap_bram_iarg_118_din1),
        .ap_bram_118_dout1(ap_bram_iarg_118_dout1),
        .ap_bram_118_we1(ap_bram_iarg_118_we1),
        .ap_bram_118_en1(ap_bram_iarg_118_en1),
        .s_axis_bram_119_tlast(s_axis_bram_119_tlast),
        .s_axis_bram_119_tvalid(s_axis_bram_119_tvalid),
        .s_axis_bram_119_tkeep(s_axis_bram_119_tkeep),
        .s_axis_bram_119_tstrb(s_axis_bram_119_tstrb),
        .s_axis_bram_119_tdata(s_axis_bram_119_tdata),
        .s_axis_bram_119_tready(s_axis_bram_119_tready),
        .ap_bram_119_addr0(ap_bram_iarg_119_addr0),
        .ap_bram_119_din0(ap_bram_iarg_119_din0),
        .ap_bram_119_dout0(ap_bram_iarg_119_dout0),
        .ap_bram_119_we0(ap_bram_iarg_119_we0),
        .ap_bram_119_en0(ap_bram_iarg_119_en0),
        .ap_bram_119_addr1(ap_bram_iarg_119_addr1),
        .ap_bram_119_din1(ap_bram_iarg_119_din1),
        .ap_bram_119_dout1(ap_bram_iarg_119_dout1),
        .ap_bram_119_we1(ap_bram_iarg_119_we1),
        .ap_bram_119_en1(ap_bram_iarg_119_en1),
        .s_axis_bram_120_tlast(s_axis_bram_120_tlast),
        .s_axis_bram_120_tvalid(s_axis_bram_120_tvalid),
        .s_axis_bram_120_tkeep(s_axis_bram_120_tkeep),
        .s_axis_bram_120_tstrb(s_axis_bram_120_tstrb),
        .s_axis_bram_120_tdata(s_axis_bram_120_tdata),
        .s_axis_bram_120_tready(s_axis_bram_120_tready),
        .ap_bram_120_addr0(ap_bram_iarg_120_addr0),
        .ap_bram_120_din0(ap_bram_iarg_120_din0),
        .ap_bram_120_dout0(ap_bram_iarg_120_dout0),
        .ap_bram_120_we0(ap_bram_iarg_120_we0),
        .ap_bram_120_en0(ap_bram_iarg_120_en0),
        .ap_bram_120_addr1(ap_bram_iarg_120_addr1),
        .ap_bram_120_din1(ap_bram_iarg_120_din1),
        .ap_bram_120_dout1(ap_bram_iarg_120_dout1),
        .ap_bram_120_we1(ap_bram_iarg_120_we1),
        .ap_bram_120_en1(ap_bram_iarg_120_en1),
        .s_axis_bram_121_tlast(s_axis_bram_121_tlast),
        .s_axis_bram_121_tvalid(s_axis_bram_121_tvalid),
        .s_axis_bram_121_tkeep(s_axis_bram_121_tkeep),
        .s_axis_bram_121_tstrb(s_axis_bram_121_tstrb),
        .s_axis_bram_121_tdata(s_axis_bram_121_tdata),
        .s_axis_bram_121_tready(s_axis_bram_121_tready),
        .ap_bram_121_addr0(ap_bram_iarg_121_addr0),
        .ap_bram_121_din0(ap_bram_iarg_121_din0),
        .ap_bram_121_dout0(ap_bram_iarg_121_dout0),
        .ap_bram_121_we0(ap_bram_iarg_121_we0),
        .ap_bram_121_en0(ap_bram_iarg_121_en0),
        .ap_bram_121_addr1(ap_bram_iarg_121_addr1),
        .ap_bram_121_din1(ap_bram_iarg_121_din1),
        .ap_bram_121_dout1(ap_bram_iarg_121_dout1),
        .ap_bram_121_we1(ap_bram_iarg_121_we1),
        .ap_bram_121_en1(ap_bram_iarg_121_en1),
        .s_axis_bram_122_tlast(s_axis_bram_122_tlast),
        .s_axis_bram_122_tvalid(s_axis_bram_122_tvalid),
        .s_axis_bram_122_tkeep(s_axis_bram_122_tkeep),
        .s_axis_bram_122_tstrb(s_axis_bram_122_tstrb),
        .s_axis_bram_122_tdata(s_axis_bram_122_tdata),
        .s_axis_bram_122_tready(s_axis_bram_122_tready),
        .ap_bram_122_addr0(ap_bram_iarg_122_addr0),
        .ap_bram_122_din0(ap_bram_iarg_122_din0),
        .ap_bram_122_dout0(ap_bram_iarg_122_dout0),
        .ap_bram_122_we0(ap_bram_iarg_122_we0),
        .ap_bram_122_en0(ap_bram_iarg_122_en0),
        .ap_bram_122_addr1(ap_bram_iarg_122_addr1),
        .ap_bram_122_din1(ap_bram_iarg_122_din1),
        .ap_bram_122_dout1(ap_bram_iarg_122_dout1),
        .ap_bram_122_we1(ap_bram_iarg_122_we1),
        .ap_bram_122_en1(ap_bram_iarg_122_en1),
        .s_axis_bram_123_tlast(s_axis_bram_123_tlast),
        .s_axis_bram_123_tvalid(s_axis_bram_123_tvalid),
        .s_axis_bram_123_tkeep(s_axis_bram_123_tkeep),
        .s_axis_bram_123_tstrb(s_axis_bram_123_tstrb),
        .s_axis_bram_123_tdata(s_axis_bram_123_tdata),
        .s_axis_bram_123_tready(s_axis_bram_123_tready),
        .ap_bram_123_addr0(ap_bram_iarg_123_addr0),
        .ap_bram_123_din0(ap_bram_iarg_123_din0),
        .ap_bram_123_dout0(ap_bram_iarg_123_dout0),
        .ap_bram_123_we0(ap_bram_iarg_123_we0),
        .ap_bram_123_en0(ap_bram_iarg_123_en0),
        .ap_bram_123_addr1(ap_bram_iarg_123_addr1),
        .ap_bram_123_din1(ap_bram_iarg_123_din1),
        .ap_bram_123_dout1(ap_bram_iarg_123_dout1),
        .ap_bram_123_we1(ap_bram_iarg_123_we1),
        .ap_bram_123_en1(ap_bram_iarg_123_en1),
        .s_axis_bram_124_tlast(s_axis_bram_124_tlast),
        .s_axis_bram_124_tvalid(s_axis_bram_124_tvalid),
        .s_axis_bram_124_tkeep(s_axis_bram_124_tkeep),
        .s_axis_bram_124_tstrb(s_axis_bram_124_tstrb),
        .s_axis_bram_124_tdata(s_axis_bram_124_tdata),
        .s_axis_bram_124_tready(s_axis_bram_124_tready),
        .ap_bram_124_addr0(ap_bram_iarg_124_addr0),
        .ap_bram_124_din0(ap_bram_iarg_124_din0),
        .ap_bram_124_dout0(ap_bram_iarg_124_dout0),
        .ap_bram_124_we0(ap_bram_iarg_124_we0),
        .ap_bram_124_en0(ap_bram_iarg_124_en0),
        .ap_bram_124_addr1(ap_bram_iarg_124_addr1),
        .ap_bram_124_din1(ap_bram_iarg_124_din1),
        .ap_bram_124_dout1(ap_bram_iarg_124_dout1),
        .ap_bram_124_we1(ap_bram_iarg_124_we1),
        .ap_bram_124_en1(ap_bram_iarg_124_en1),
        .s_axis_bram_125_tlast(s_axis_bram_125_tlast),
        .s_axis_bram_125_tvalid(s_axis_bram_125_tvalid),
        .s_axis_bram_125_tkeep(s_axis_bram_125_tkeep),
        .s_axis_bram_125_tstrb(s_axis_bram_125_tstrb),
        .s_axis_bram_125_tdata(s_axis_bram_125_tdata),
        .s_axis_bram_125_tready(s_axis_bram_125_tready),
        .ap_bram_125_addr0(ap_bram_iarg_125_addr0),
        .ap_bram_125_din0(ap_bram_iarg_125_din0),
        .ap_bram_125_dout0(ap_bram_iarg_125_dout0),
        .ap_bram_125_we0(ap_bram_iarg_125_we0),
        .ap_bram_125_en0(ap_bram_iarg_125_en0),
        .ap_bram_125_addr1(ap_bram_iarg_125_addr1),
        .ap_bram_125_din1(ap_bram_iarg_125_din1),
        .ap_bram_125_dout1(ap_bram_iarg_125_dout1),
        .ap_bram_125_we1(ap_bram_iarg_125_we1),
        .ap_bram_125_en1(ap_bram_iarg_125_en1),
        .s_axis_bram_126_tlast(s_axis_bram_126_tlast),
        .s_axis_bram_126_tvalid(s_axis_bram_126_tvalid),
        .s_axis_bram_126_tkeep(s_axis_bram_126_tkeep),
        .s_axis_bram_126_tstrb(s_axis_bram_126_tstrb),
        .s_axis_bram_126_tdata(s_axis_bram_126_tdata),
        .s_axis_bram_126_tready(s_axis_bram_126_tready),
        .ap_bram_126_addr0(ap_bram_iarg_126_addr0),
        .ap_bram_126_din0(ap_bram_iarg_126_din0),
        .ap_bram_126_dout0(ap_bram_iarg_126_dout0),
        .ap_bram_126_we0(ap_bram_iarg_126_we0),
        .ap_bram_126_en0(ap_bram_iarg_126_en0),
        .ap_bram_126_addr1(ap_bram_iarg_126_addr1),
        .ap_bram_126_din1(ap_bram_iarg_126_din1),
        .ap_bram_126_dout1(ap_bram_iarg_126_dout1),
        .ap_bram_126_we1(ap_bram_iarg_126_we1),
        .ap_bram_126_en1(ap_bram_iarg_126_en1),
        .s_axis_bram_127_tlast(s_axis_bram_127_tlast),
        .s_axis_bram_127_tvalid(s_axis_bram_127_tvalid),
        .s_axis_bram_127_tkeep(s_axis_bram_127_tkeep),
        .s_axis_bram_127_tstrb(s_axis_bram_127_tstrb),
        .s_axis_bram_127_tdata(s_axis_bram_127_tdata),
        .s_axis_bram_127_tready(s_axis_bram_127_tready),
        .ap_bram_127_addr0(ap_bram_iarg_127_addr0),
        .ap_bram_127_din0(ap_bram_iarg_127_din0),
        .ap_bram_127_dout0(ap_bram_iarg_127_dout0),
        .ap_bram_127_we0(ap_bram_iarg_127_we0),
        .ap_bram_127_en0(ap_bram_iarg_127_en0),
        .ap_bram_127_addr1(ap_bram_iarg_127_addr1),
        .ap_bram_127_din1(ap_bram_iarg_127_din1),
        .ap_bram_127_dout1(ap_bram_iarg_127_dout1),
        .ap_bram_127_we1(ap_bram_iarg_127_we1),
        .ap_bram_127_en1(ap_bram_iarg_127_en1),
        .m_axis_bram_0_tlast(m_axis_bramio_0_tlast),
        .m_axis_bram_0_tvalid(m_axis_bramio_0_tvalid),
        .m_axis_bram_0_tkeep(m_axis_bramio_0_tkeep),
        .m_axis_bram_0_tstrb(m_axis_bramio_0_tstrb),
        .m_axis_bram_0_tdata(m_axis_bramio_0_tdata),
        .m_axis_bram_0_tready(m_axis_bramio_0_tready),
        .m_axis_bram_1_tlast(m_axis_bramio_1_tlast),
        .m_axis_bram_1_tvalid(m_axis_bramio_1_tvalid),
        .m_axis_bram_1_tkeep(m_axis_bramio_1_tkeep),
        .m_axis_bram_1_tstrb(m_axis_bramio_1_tstrb),
        .m_axis_bram_1_tdata(m_axis_bramio_1_tdata),
        .m_axis_bram_1_tready(m_axis_bramio_1_tready),
        .m_axis_bram_2_tlast(m_axis_bramio_2_tlast),
        .m_axis_bram_2_tvalid(m_axis_bramio_2_tvalid),
        .m_axis_bram_2_tkeep(m_axis_bramio_2_tkeep),
        .m_axis_bram_2_tstrb(m_axis_bramio_2_tstrb),
        .m_axis_bram_2_tdata(m_axis_bramio_2_tdata),
        .m_axis_bram_2_tready(m_axis_bramio_2_tready),
        .m_axis_bram_3_tlast(m_axis_bramio_3_tlast),
        .m_axis_bram_3_tvalid(m_axis_bramio_3_tvalid),
        .m_axis_bram_3_tkeep(m_axis_bramio_3_tkeep),
        .m_axis_bram_3_tstrb(m_axis_bramio_3_tstrb),
        .m_axis_bram_3_tdata(m_axis_bramio_3_tdata),
        .m_axis_bram_3_tready(m_axis_bramio_3_tready),
        .m_axis_bram_4_tlast(m_axis_bramio_4_tlast),
        .m_axis_bram_4_tvalid(m_axis_bramio_4_tvalid),
        .m_axis_bram_4_tkeep(m_axis_bramio_4_tkeep),
        .m_axis_bram_4_tstrb(m_axis_bramio_4_tstrb),
        .m_axis_bram_4_tdata(m_axis_bramio_4_tdata),
        .m_axis_bram_4_tready(m_axis_bramio_4_tready),
        .m_axis_bram_5_tlast(m_axis_bramio_5_tlast),
        .m_axis_bram_5_tvalid(m_axis_bramio_5_tvalid),
        .m_axis_bram_5_tkeep(m_axis_bramio_5_tkeep),
        .m_axis_bram_5_tstrb(m_axis_bramio_5_tstrb),
        .m_axis_bram_5_tdata(m_axis_bramio_5_tdata),
        .m_axis_bram_5_tready(m_axis_bramio_5_tready),
        .m_axis_bram_6_tlast(m_axis_bramio_6_tlast),
        .m_axis_bram_6_tvalid(m_axis_bramio_6_tvalid),
        .m_axis_bram_6_tkeep(m_axis_bramio_6_tkeep),
        .m_axis_bram_6_tstrb(m_axis_bramio_6_tstrb),
        .m_axis_bram_6_tdata(m_axis_bramio_6_tdata),
        .m_axis_bram_6_tready(m_axis_bramio_6_tready),
        .m_axis_bram_7_tlast(m_axis_bramio_7_tlast),
        .m_axis_bram_7_tvalid(m_axis_bramio_7_tvalid),
        .m_axis_bram_7_tkeep(m_axis_bramio_7_tkeep),
        .m_axis_bram_7_tstrb(m_axis_bramio_7_tstrb),
        .m_axis_bram_7_tdata(m_axis_bramio_7_tdata),
        .m_axis_bram_7_tready(m_axis_bramio_7_tready),
        .m_axis_bram_8_tlast(m_axis_bramio_8_tlast),
        .m_axis_bram_8_tvalid(m_axis_bramio_8_tvalid),
        .m_axis_bram_8_tkeep(m_axis_bramio_8_tkeep),
        .m_axis_bram_8_tstrb(m_axis_bramio_8_tstrb),
        .m_axis_bram_8_tdata(m_axis_bramio_8_tdata),
        .m_axis_bram_8_tready(m_axis_bramio_8_tready),
        .m_axis_bram_9_tlast(m_axis_bramio_9_tlast),
        .m_axis_bram_9_tvalid(m_axis_bramio_9_tvalid),
        .m_axis_bram_9_tkeep(m_axis_bramio_9_tkeep),
        .m_axis_bram_9_tstrb(m_axis_bramio_9_tstrb),
        .m_axis_bram_9_tdata(m_axis_bramio_9_tdata),
        .m_axis_bram_9_tready(m_axis_bramio_9_tready),
        .m_axis_bram_10_tlast(m_axis_bramio_10_tlast),
        .m_axis_bram_10_tvalid(m_axis_bramio_10_tvalid),
        .m_axis_bram_10_tkeep(m_axis_bramio_10_tkeep),
        .m_axis_bram_10_tstrb(m_axis_bramio_10_tstrb),
        .m_axis_bram_10_tdata(m_axis_bramio_10_tdata),
        .m_axis_bram_10_tready(m_axis_bramio_10_tready),
        .m_axis_bram_11_tlast(m_axis_bramio_11_tlast),
        .m_axis_bram_11_tvalid(m_axis_bramio_11_tvalid),
        .m_axis_bram_11_tkeep(m_axis_bramio_11_tkeep),
        .m_axis_bram_11_tstrb(m_axis_bramio_11_tstrb),
        .m_axis_bram_11_tdata(m_axis_bramio_11_tdata),
        .m_axis_bram_11_tready(m_axis_bramio_11_tready),
        .m_axis_bram_12_tlast(m_axis_bramio_12_tlast),
        .m_axis_bram_12_tvalid(m_axis_bramio_12_tvalid),
        .m_axis_bram_12_tkeep(m_axis_bramio_12_tkeep),
        .m_axis_bram_12_tstrb(m_axis_bramio_12_tstrb),
        .m_axis_bram_12_tdata(m_axis_bramio_12_tdata),
        .m_axis_bram_12_tready(m_axis_bramio_12_tready),
        .m_axis_bram_13_tlast(m_axis_bramio_13_tlast),
        .m_axis_bram_13_tvalid(m_axis_bramio_13_tvalid),
        .m_axis_bram_13_tkeep(m_axis_bramio_13_tkeep),
        .m_axis_bram_13_tstrb(m_axis_bramio_13_tstrb),
        .m_axis_bram_13_tdata(m_axis_bramio_13_tdata),
        .m_axis_bram_13_tready(m_axis_bramio_13_tready),
        .m_axis_bram_14_tlast(m_axis_bramio_14_tlast),
        .m_axis_bram_14_tvalid(m_axis_bramio_14_tvalid),
        .m_axis_bram_14_tkeep(m_axis_bramio_14_tkeep),
        .m_axis_bram_14_tstrb(m_axis_bramio_14_tstrb),
        .m_axis_bram_14_tdata(m_axis_bramio_14_tdata),
        .m_axis_bram_14_tready(m_axis_bramio_14_tready),
        .m_axis_bram_15_tlast(m_axis_bramio_15_tlast),
        .m_axis_bram_15_tvalid(m_axis_bramio_15_tvalid),
        .m_axis_bram_15_tkeep(m_axis_bramio_15_tkeep),
        .m_axis_bram_15_tstrb(m_axis_bramio_15_tstrb),
        .m_axis_bram_15_tdata(m_axis_bramio_15_tdata),
        .m_axis_bram_15_tready(m_axis_bramio_15_tready),
        .m_axis_bram_16_tlast(m_axis_bramio_16_tlast),
        .m_axis_bram_16_tvalid(m_axis_bramio_16_tvalid),
        .m_axis_bram_16_tkeep(m_axis_bramio_16_tkeep),
        .m_axis_bram_16_tstrb(m_axis_bramio_16_tstrb),
        .m_axis_bram_16_tdata(m_axis_bramio_16_tdata),
        .m_axis_bram_16_tready(m_axis_bramio_16_tready),
        .m_axis_bram_17_tlast(m_axis_bramio_17_tlast),
        .m_axis_bram_17_tvalid(m_axis_bramio_17_tvalid),
        .m_axis_bram_17_tkeep(m_axis_bramio_17_tkeep),
        .m_axis_bram_17_tstrb(m_axis_bramio_17_tstrb),
        .m_axis_bram_17_tdata(m_axis_bramio_17_tdata),
        .m_axis_bram_17_tready(m_axis_bramio_17_tready),
        .m_axis_bram_18_tlast(m_axis_bramio_18_tlast),
        .m_axis_bram_18_tvalid(m_axis_bramio_18_tvalid),
        .m_axis_bram_18_tkeep(m_axis_bramio_18_tkeep),
        .m_axis_bram_18_tstrb(m_axis_bramio_18_tstrb),
        .m_axis_bram_18_tdata(m_axis_bramio_18_tdata),
        .m_axis_bram_18_tready(m_axis_bramio_18_tready),
        .m_axis_bram_19_tlast(m_axis_bramio_19_tlast),
        .m_axis_bram_19_tvalid(m_axis_bramio_19_tvalid),
        .m_axis_bram_19_tkeep(m_axis_bramio_19_tkeep),
        .m_axis_bram_19_tstrb(m_axis_bramio_19_tstrb),
        .m_axis_bram_19_tdata(m_axis_bramio_19_tdata),
        .m_axis_bram_19_tready(m_axis_bramio_19_tready),
        .m_axis_bram_20_tlast(m_axis_bramio_20_tlast),
        .m_axis_bram_20_tvalid(m_axis_bramio_20_tvalid),
        .m_axis_bram_20_tkeep(m_axis_bramio_20_tkeep),
        .m_axis_bram_20_tstrb(m_axis_bramio_20_tstrb),
        .m_axis_bram_20_tdata(m_axis_bramio_20_tdata),
        .m_axis_bram_20_tready(m_axis_bramio_20_tready),
        .m_axis_bram_21_tlast(m_axis_bramio_21_tlast),
        .m_axis_bram_21_tvalid(m_axis_bramio_21_tvalid),
        .m_axis_bram_21_tkeep(m_axis_bramio_21_tkeep),
        .m_axis_bram_21_tstrb(m_axis_bramio_21_tstrb),
        .m_axis_bram_21_tdata(m_axis_bramio_21_tdata),
        .m_axis_bram_21_tready(m_axis_bramio_21_tready),
        .m_axis_bram_22_tlast(m_axis_bramio_22_tlast),
        .m_axis_bram_22_tvalid(m_axis_bramio_22_tvalid),
        .m_axis_bram_22_tkeep(m_axis_bramio_22_tkeep),
        .m_axis_bram_22_tstrb(m_axis_bramio_22_tstrb),
        .m_axis_bram_22_tdata(m_axis_bramio_22_tdata),
        .m_axis_bram_22_tready(m_axis_bramio_22_tready),
        .m_axis_bram_23_tlast(m_axis_bramio_23_tlast),
        .m_axis_bram_23_tvalid(m_axis_bramio_23_tvalid),
        .m_axis_bram_23_tkeep(m_axis_bramio_23_tkeep),
        .m_axis_bram_23_tstrb(m_axis_bramio_23_tstrb),
        .m_axis_bram_23_tdata(m_axis_bramio_23_tdata),
        .m_axis_bram_23_tready(m_axis_bramio_23_tready),
        .m_axis_bram_24_tlast(m_axis_bramio_24_tlast),
        .m_axis_bram_24_tvalid(m_axis_bramio_24_tvalid),
        .m_axis_bram_24_tkeep(m_axis_bramio_24_tkeep),
        .m_axis_bram_24_tstrb(m_axis_bramio_24_tstrb),
        .m_axis_bram_24_tdata(m_axis_bramio_24_tdata),
        .m_axis_bram_24_tready(m_axis_bramio_24_tready),
        .m_axis_bram_25_tlast(m_axis_bramio_25_tlast),
        .m_axis_bram_25_tvalid(m_axis_bramio_25_tvalid),
        .m_axis_bram_25_tkeep(m_axis_bramio_25_tkeep),
        .m_axis_bram_25_tstrb(m_axis_bramio_25_tstrb),
        .m_axis_bram_25_tdata(m_axis_bramio_25_tdata),
        .m_axis_bram_25_tready(m_axis_bramio_25_tready),
        .m_axis_bram_26_tlast(m_axis_bramio_26_tlast),
        .m_axis_bram_26_tvalid(m_axis_bramio_26_tvalid),
        .m_axis_bram_26_tkeep(m_axis_bramio_26_tkeep),
        .m_axis_bram_26_tstrb(m_axis_bramio_26_tstrb),
        .m_axis_bram_26_tdata(m_axis_bramio_26_tdata),
        .m_axis_bram_26_tready(m_axis_bramio_26_tready),
        .m_axis_bram_27_tlast(m_axis_bramio_27_tlast),
        .m_axis_bram_27_tvalid(m_axis_bramio_27_tvalid),
        .m_axis_bram_27_tkeep(m_axis_bramio_27_tkeep),
        .m_axis_bram_27_tstrb(m_axis_bramio_27_tstrb),
        .m_axis_bram_27_tdata(m_axis_bramio_27_tdata),
        .m_axis_bram_27_tready(m_axis_bramio_27_tready),
        .m_axis_bram_28_tlast(m_axis_bramio_28_tlast),
        .m_axis_bram_28_tvalid(m_axis_bramio_28_tvalid),
        .m_axis_bram_28_tkeep(m_axis_bramio_28_tkeep),
        .m_axis_bram_28_tstrb(m_axis_bramio_28_tstrb),
        .m_axis_bram_28_tdata(m_axis_bramio_28_tdata),
        .m_axis_bram_28_tready(m_axis_bramio_28_tready),
        .m_axis_bram_29_tlast(m_axis_bramio_29_tlast),
        .m_axis_bram_29_tvalid(m_axis_bramio_29_tvalid),
        .m_axis_bram_29_tkeep(m_axis_bramio_29_tkeep),
        .m_axis_bram_29_tstrb(m_axis_bramio_29_tstrb),
        .m_axis_bram_29_tdata(m_axis_bramio_29_tdata),
        .m_axis_bram_29_tready(m_axis_bramio_29_tready),
        .m_axis_bram_30_tlast(m_axis_bramio_30_tlast),
        .m_axis_bram_30_tvalid(m_axis_bramio_30_tvalid),
        .m_axis_bram_30_tkeep(m_axis_bramio_30_tkeep),
        .m_axis_bram_30_tstrb(m_axis_bramio_30_tstrb),
        .m_axis_bram_30_tdata(m_axis_bramio_30_tdata),
        .m_axis_bram_30_tready(m_axis_bramio_30_tready),
        .m_axis_bram_31_tlast(m_axis_bramio_31_tlast),
        .m_axis_bram_31_tvalid(m_axis_bramio_31_tvalid),
        .m_axis_bram_31_tkeep(m_axis_bramio_31_tkeep),
        .m_axis_bram_31_tstrb(m_axis_bramio_31_tstrb),
        .m_axis_bram_31_tdata(m_axis_bramio_31_tdata),
        .m_axis_bram_31_tready(m_axis_bramio_31_tready),
        .m_axis_bram_32_tlast(m_axis_bramio_32_tlast),
        .m_axis_bram_32_tvalid(m_axis_bramio_32_tvalid),
        .m_axis_bram_32_tkeep(m_axis_bramio_32_tkeep),
        .m_axis_bram_32_tstrb(m_axis_bramio_32_tstrb),
        .m_axis_bram_32_tdata(m_axis_bramio_32_tdata),
        .m_axis_bram_32_tready(m_axis_bramio_32_tready),
        .m_axis_bram_33_tlast(m_axis_bramio_33_tlast),
        .m_axis_bram_33_tvalid(m_axis_bramio_33_tvalid),
        .m_axis_bram_33_tkeep(m_axis_bramio_33_tkeep),
        .m_axis_bram_33_tstrb(m_axis_bramio_33_tstrb),
        .m_axis_bram_33_tdata(m_axis_bramio_33_tdata),
        .m_axis_bram_33_tready(m_axis_bramio_33_tready),
        .m_axis_bram_34_tlast(m_axis_bramio_34_tlast),
        .m_axis_bram_34_tvalid(m_axis_bramio_34_tvalid),
        .m_axis_bram_34_tkeep(m_axis_bramio_34_tkeep),
        .m_axis_bram_34_tstrb(m_axis_bramio_34_tstrb),
        .m_axis_bram_34_tdata(m_axis_bramio_34_tdata),
        .m_axis_bram_34_tready(m_axis_bramio_34_tready),
        .m_axis_bram_35_tlast(m_axis_bramio_35_tlast),
        .m_axis_bram_35_tvalid(m_axis_bramio_35_tvalid),
        .m_axis_bram_35_tkeep(m_axis_bramio_35_tkeep),
        .m_axis_bram_35_tstrb(m_axis_bramio_35_tstrb),
        .m_axis_bram_35_tdata(m_axis_bramio_35_tdata),
        .m_axis_bram_35_tready(m_axis_bramio_35_tready),
        .m_axis_bram_36_tlast(m_axis_bramio_36_tlast),
        .m_axis_bram_36_tvalid(m_axis_bramio_36_tvalid),
        .m_axis_bram_36_tkeep(m_axis_bramio_36_tkeep),
        .m_axis_bram_36_tstrb(m_axis_bramio_36_tstrb),
        .m_axis_bram_36_tdata(m_axis_bramio_36_tdata),
        .m_axis_bram_36_tready(m_axis_bramio_36_tready),
        .m_axis_bram_37_tlast(m_axis_bramio_37_tlast),
        .m_axis_bram_37_tvalid(m_axis_bramio_37_tvalid),
        .m_axis_bram_37_tkeep(m_axis_bramio_37_tkeep),
        .m_axis_bram_37_tstrb(m_axis_bramio_37_tstrb),
        .m_axis_bram_37_tdata(m_axis_bramio_37_tdata),
        .m_axis_bram_37_tready(m_axis_bramio_37_tready),
        .m_axis_bram_38_tlast(m_axis_bramio_38_tlast),
        .m_axis_bram_38_tvalid(m_axis_bramio_38_tvalid),
        .m_axis_bram_38_tkeep(m_axis_bramio_38_tkeep),
        .m_axis_bram_38_tstrb(m_axis_bramio_38_tstrb),
        .m_axis_bram_38_tdata(m_axis_bramio_38_tdata),
        .m_axis_bram_38_tready(m_axis_bramio_38_tready),
        .m_axis_bram_39_tlast(m_axis_bramio_39_tlast),
        .m_axis_bram_39_tvalid(m_axis_bramio_39_tvalid),
        .m_axis_bram_39_tkeep(m_axis_bramio_39_tkeep),
        .m_axis_bram_39_tstrb(m_axis_bramio_39_tstrb),
        .m_axis_bram_39_tdata(m_axis_bramio_39_tdata),
        .m_axis_bram_39_tready(m_axis_bramio_39_tready),
        .m_axis_bram_40_tlast(m_axis_bramio_40_tlast),
        .m_axis_bram_40_tvalid(m_axis_bramio_40_tvalid),
        .m_axis_bram_40_tkeep(m_axis_bramio_40_tkeep),
        .m_axis_bram_40_tstrb(m_axis_bramio_40_tstrb),
        .m_axis_bram_40_tdata(m_axis_bramio_40_tdata),
        .m_axis_bram_40_tready(m_axis_bramio_40_tready),
        .m_axis_bram_41_tlast(m_axis_bramio_41_tlast),
        .m_axis_bram_41_tvalid(m_axis_bramio_41_tvalid),
        .m_axis_bram_41_tkeep(m_axis_bramio_41_tkeep),
        .m_axis_bram_41_tstrb(m_axis_bramio_41_tstrb),
        .m_axis_bram_41_tdata(m_axis_bramio_41_tdata),
        .m_axis_bram_41_tready(m_axis_bramio_41_tready),
        .m_axis_bram_42_tlast(m_axis_bramio_42_tlast),
        .m_axis_bram_42_tvalid(m_axis_bramio_42_tvalid),
        .m_axis_bram_42_tkeep(m_axis_bramio_42_tkeep),
        .m_axis_bram_42_tstrb(m_axis_bramio_42_tstrb),
        .m_axis_bram_42_tdata(m_axis_bramio_42_tdata),
        .m_axis_bram_42_tready(m_axis_bramio_42_tready),
        .m_axis_bram_43_tlast(m_axis_bramio_43_tlast),
        .m_axis_bram_43_tvalid(m_axis_bramio_43_tvalid),
        .m_axis_bram_43_tkeep(m_axis_bramio_43_tkeep),
        .m_axis_bram_43_tstrb(m_axis_bramio_43_tstrb),
        .m_axis_bram_43_tdata(m_axis_bramio_43_tdata),
        .m_axis_bram_43_tready(m_axis_bramio_43_tready),
        .m_axis_bram_44_tlast(m_axis_bramio_44_tlast),
        .m_axis_bram_44_tvalid(m_axis_bramio_44_tvalid),
        .m_axis_bram_44_tkeep(m_axis_bramio_44_tkeep),
        .m_axis_bram_44_tstrb(m_axis_bramio_44_tstrb),
        .m_axis_bram_44_tdata(m_axis_bramio_44_tdata),
        .m_axis_bram_44_tready(m_axis_bramio_44_tready),
        .m_axis_bram_45_tlast(m_axis_bramio_45_tlast),
        .m_axis_bram_45_tvalid(m_axis_bramio_45_tvalid),
        .m_axis_bram_45_tkeep(m_axis_bramio_45_tkeep),
        .m_axis_bram_45_tstrb(m_axis_bramio_45_tstrb),
        .m_axis_bram_45_tdata(m_axis_bramio_45_tdata),
        .m_axis_bram_45_tready(m_axis_bramio_45_tready),
        .m_axis_bram_46_tlast(m_axis_bramio_46_tlast),
        .m_axis_bram_46_tvalid(m_axis_bramio_46_tvalid),
        .m_axis_bram_46_tkeep(m_axis_bramio_46_tkeep),
        .m_axis_bram_46_tstrb(m_axis_bramio_46_tstrb),
        .m_axis_bram_46_tdata(m_axis_bramio_46_tdata),
        .m_axis_bram_46_tready(m_axis_bramio_46_tready),
        .m_axis_bram_47_tlast(m_axis_bramio_47_tlast),
        .m_axis_bram_47_tvalid(m_axis_bramio_47_tvalid),
        .m_axis_bram_47_tkeep(m_axis_bramio_47_tkeep),
        .m_axis_bram_47_tstrb(m_axis_bramio_47_tstrb),
        .m_axis_bram_47_tdata(m_axis_bramio_47_tdata),
        .m_axis_bram_47_tready(m_axis_bramio_47_tready),
        .m_axis_bram_48_tlast(m_axis_bramio_48_tlast),
        .m_axis_bram_48_tvalid(m_axis_bramio_48_tvalid),
        .m_axis_bram_48_tkeep(m_axis_bramio_48_tkeep),
        .m_axis_bram_48_tstrb(m_axis_bramio_48_tstrb),
        .m_axis_bram_48_tdata(m_axis_bramio_48_tdata),
        .m_axis_bram_48_tready(m_axis_bramio_48_tready),
        .m_axis_bram_49_tlast(m_axis_bramio_49_tlast),
        .m_axis_bram_49_tvalid(m_axis_bramio_49_tvalid),
        .m_axis_bram_49_tkeep(m_axis_bramio_49_tkeep),
        .m_axis_bram_49_tstrb(m_axis_bramio_49_tstrb),
        .m_axis_bram_49_tdata(m_axis_bramio_49_tdata),
        .m_axis_bram_49_tready(m_axis_bramio_49_tready),
        .m_axis_bram_50_tlast(m_axis_bramio_50_tlast),
        .m_axis_bram_50_tvalid(m_axis_bramio_50_tvalid),
        .m_axis_bram_50_tkeep(m_axis_bramio_50_tkeep),
        .m_axis_bram_50_tstrb(m_axis_bramio_50_tstrb),
        .m_axis_bram_50_tdata(m_axis_bramio_50_tdata),
        .m_axis_bram_50_tready(m_axis_bramio_50_tready),
        .m_axis_bram_51_tlast(m_axis_bramio_51_tlast),
        .m_axis_bram_51_tvalid(m_axis_bramio_51_tvalid),
        .m_axis_bram_51_tkeep(m_axis_bramio_51_tkeep),
        .m_axis_bram_51_tstrb(m_axis_bramio_51_tstrb),
        .m_axis_bram_51_tdata(m_axis_bramio_51_tdata),
        .m_axis_bram_51_tready(m_axis_bramio_51_tready),
        .m_axis_bram_52_tlast(m_axis_bramio_52_tlast),
        .m_axis_bram_52_tvalid(m_axis_bramio_52_tvalid),
        .m_axis_bram_52_tkeep(m_axis_bramio_52_tkeep),
        .m_axis_bram_52_tstrb(m_axis_bramio_52_tstrb),
        .m_axis_bram_52_tdata(m_axis_bramio_52_tdata),
        .m_axis_bram_52_tready(m_axis_bramio_52_tready),
        .m_axis_bram_53_tlast(m_axis_bramio_53_tlast),
        .m_axis_bram_53_tvalid(m_axis_bramio_53_tvalid),
        .m_axis_bram_53_tkeep(m_axis_bramio_53_tkeep),
        .m_axis_bram_53_tstrb(m_axis_bramio_53_tstrb),
        .m_axis_bram_53_tdata(m_axis_bramio_53_tdata),
        .m_axis_bram_53_tready(m_axis_bramio_53_tready),
        .m_axis_bram_54_tlast(m_axis_bramio_54_tlast),
        .m_axis_bram_54_tvalid(m_axis_bramio_54_tvalid),
        .m_axis_bram_54_tkeep(m_axis_bramio_54_tkeep),
        .m_axis_bram_54_tstrb(m_axis_bramio_54_tstrb),
        .m_axis_bram_54_tdata(m_axis_bramio_54_tdata),
        .m_axis_bram_54_tready(m_axis_bramio_54_tready),
        .m_axis_bram_55_tlast(m_axis_bramio_55_tlast),
        .m_axis_bram_55_tvalid(m_axis_bramio_55_tvalid),
        .m_axis_bram_55_tkeep(m_axis_bramio_55_tkeep),
        .m_axis_bram_55_tstrb(m_axis_bramio_55_tstrb),
        .m_axis_bram_55_tdata(m_axis_bramio_55_tdata),
        .m_axis_bram_55_tready(m_axis_bramio_55_tready),
        .m_axis_bram_56_tlast(m_axis_bramio_56_tlast),
        .m_axis_bram_56_tvalid(m_axis_bramio_56_tvalid),
        .m_axis_bram_56_tkeep(m_axis_bramio_56_tkeep),
        .m_axis_bram_56_tstrb(m_axis_bramio_56_tstrb),
        .m_axis_bram_56_tdata(m_axis_bramio_56_tdata),
        .m_axis_bram_56_tready(m_axis_bramio_56_tready),
        .m_axis_bram_57_tlast(m_axis_bramio_57_tlast),
        .m_axis_bram_57_tvalid(m_axis_bramio_57_tvalid),
        .m_axis_bram_57_tkeep(m_axis_bramio_57_tkeep),
        .m_axis_bram_57_tstrb(m_axis_bramio_57_tstrb),
        .m_axis_bram_57_tdata(m_axis_bramio_57_tdata),
        .m_axis_bram_57_tready(m_axis_bramio_57_tready),
        .m_axis_bram_58_tlast(m_axis_bramio_58_tlast),
        .m_axis_bram_58_tvalid(m_axis_bramio_58_tvalid),
        .m_axis_bram_58_tkeep(m_axis_bramio_58_tkeep),
        .m_axis_bram_58_tstrb(m_axis_bramio_58_tstrb),
        .m_axis_bram_58_tdata(m_axis_bramio_58_tdata),
        .m_axis_bram_58_tready(m_axis_bramio_58_tready),
        .m_axis_bram_59_tlast(m_axis_bramio_59_tlast),
        .m_axis_bram_59_tvalid(m_axis_bramio_59_tvalid),
        .m_axis_bram_59_tkeep(m_axis_bramio_59_tkeep),
        .m_axis_bram_59_tstrb(m_axis_bramio_59_tstrb),
        .m_axis_bram_59_tdata(m_axis_bramio_59_tdata),
        .m_axis_bram_59_tready(m_axis_bramio_59_tready),
        .m_axis_bram_60_tlast(m_axis_bramio_60_tlast),
        .m_axis_bram_60_tvalid(m_axis_bramio_60_tvalid),
        .m_axis_bram_60_tkeep(m_axis_bramio_60_tkeep),
        .m_axis_bram_60_tstrb(m_axis_bramio_60_tstrb),
        .m_axis_bram_60_tdata(m_axis_bramio_60_tdata),
        .m_axis_bram_60_tready(m_axis_bramio_60_tready),
        .m_axis_bram_61_tlast(m_axis_bramio_61_tlast),
        .m_axis_bram_61_tvalid(m_axis_bramio_61_tvalid),
        .m_axis_bram_61_tkeep(m_axis_bramio_61_tkeep),
        .m_axis_bram_61_tstrb(m_axis_bramio_61_tstrb),
        .m_axis_bram_61_tdata(m_axis_bramio_61_tdata),
        .m_axis_bram_61_tready(m_axis_bramio_61_tready),
        .m_axis_bram_62_tlast(m_axis_bramio_62_tlast),
        .m_axis_bram_62_tvalid(m_axis_bramio_62_tvalid),
        .m_axis_bram_62_tkeep(m_axis_bramio_62_tkeep),
        .m_axis_bram_62_tstrb(m_axis_bramio_62_tstrb),
        .m_axis_bram_62_tdata(m_axis_bramio_62_tdata),
        .m_axis_bram_62_tready(m_axis_bramio_62_tready),
        .m_axis_bram_63_tlast(m_axis_bramio_63_tlast),
        .m_axis_bram_63_tvalid(m_axis_bramio_63_tvalid),
        .m_axis_bram_63_tkeep(m_axis_bramio_63_tkeep),
        .m_axis_bram_63_tstrb(m_axis_bramio_63_tstrb),
        .m_axis_bram_63_tdata(m_axis_bramio_63_tdata),
        .m_axis_bram_63_tready(m_axis_bramio_63_tready),
        .m_axis_bram_64_tlast(m_axis_bramio_64_tlast),
        .m_axis_bram_64_tvalid(m_axis_bramio_64_tvalid),
        .m_axis_bram_64_tkeep(m_axis_bramio_64_tkeep),
        .m_axis_bram_64_tstrb(m_axis_bramio_64_tstrb),
        .m_axis_bram_64_tdata(m_axis_bramio_64_tdata),
        .m_axis_bram_64_tready(m_axis_bramio_64_tready),
        .m_axis_bram_65_tlast(m_axis_bramio_65_tlast),
        .m_axis_bram_65_tvalid(m_axis_bramio_65_tvalid),
        .m_axis_bram_65_tkeep(m_axis_bramio_65_tkeep),
        .m_axis_bram_65_tstrb(m_axis_bramio_65_tstrb),
        .m_axis_bram_65_tdata(m_axis_bramio_65_tdata),
        .m_axis_bram_65_tready(m_axis_bramio_65_tready),
        .m_axis_bram_66_tlast(m_axis_bramio_66_tlast),
        .m_axis_bram_66_tvalid(m_axis_bramio_66_tvalid),
        .m_axis_bram_66_tkeep(m_axis_bramio_66_tkeep),
        .m_axis_bram_66_tstrb(m_axis_bramio_66_tstrb),
        .m_axis_bram_66_tdata(m_axis_bramio_66_tdata),
        .m_axis_bram_66_tready(m_axis_bramio_66_tready),
        .m_axis_bram_67_tlast(m_axis_bramio_67_tlast),
        .m_axis_bram_67_tvalid(m_axis_bramio_67_tvalid),
        .m_axis_bram_67_tkeep(m_axis_bramio_67_tkeep),
        .m_axis_bram_67_tstrb(m_axis_bramio_67_tstrb),
        .m_axis_bram_67_tdata(m_axis_bramio_67_tdata),
        .m_axis_bram_67_tready(m_axis_bramio_67_tready),
        .m_axis_bram_68_tlast(m_axis_bramio_68_tlast),
        .m_axis_bram_68_tvalid(m_axis_bramio_68_tvalid),
        .m_axis_bram_68_tkeep(m_axis_bramio_68_tkeep),
        .m_axis_bram_68_tstrb(m_axis_bramio_68_tstrb),
        .m_axis_bram_68_tdata(m_axis_bramio_68_tdata),
        .m_axis_bram_68_tready(m_axis_bramio_68_tready),
        .m_axis_bram_69_tlast(m_axis_bramio_69_tlast),
        .m_axis_bram_69_tvalid(m_axis_bramio_69_tvalid),
        .m_axis_bram_69_tkeep(m_axis_bramio_69_tkeep),
        .m_axis_bram_69_tstrb(m_axis_bramio_69_tstrb),
        .m_axis_bram_69_tdata(m_axis_bramio_69_tdata),
        .m_axis_bram_69_tready(m_axis_bramio_69_tready),
        .m_axis_bram_70_tlast(m_axis_bramio_70_tlast),
        .m_axis_bram_70_tvalid(m_axis_bramio_70_tvalid),
        .m_axis_bram_70_tkeep(m_axis_bramio_70_tkeep),
        .m_axis_bram_70_tstrb(m_axis_bramio_70_tstrb),
        .m_axis_bram_70_tdata(m_axis_bramio_70_tdata),
        .m_axis_bram_70_tready(m_axis_bramio_70_tready),
        .m_axis_bram_71_tlast(m_axis_bramio_71_tlast),
        .m_axis_bram_71_tvalid(m_axis_bramio_71_tvalid),
        .m_axis_bram_71_tkeep(m_axis_bramio_71_tkeep),
        .m_axis_bram_71_tstrb(m_axis_bramio_71_tstrb),
        .m_axis_bram_71_tdata(m_axis_bramio_71_tdata),
        .m_axis_bram_71_tready(m_axis_bramio_71_tready),
        .m_axis_bram_72_tlast(m_axis_bramio_72_tlast),
        .m_axis_bram_72_tvalid(m_axis_bramio_72_tvalid),
        .m_axis_bram_72_tkeep(m_axis_bramio_72_tkeep),
        .m_axis_bram_72_tstrb(m_axis_bramio_72_tstrb),
        .m_axis_bram_72_tdata(m_axis_bramio_72_tdata),
        .m_axis_bram_72_tready(m_axis_bramio_72_tready),
        .m_axis_bram_73_tlast(m_axis_bramio_73_tlast),
        .m_axis_bram_73_tvalid(m_axis_bramio_73_tvalid),
        .m_axis_bram_73_tkeep(m_axis_bramio_73_tkeep),
        .m_axis_bram_73_tstrb(m_axis_bramio_73_tstrb),
        .m_axis_bram_73_tdata(m_axis_bramio_73_tdata),
        .m_axis_bram_73_tready(m_axis_bramio_73_tready),
        .m_axis_bram_74_tlast(m_axis_bramio_74_tlast),
        .m_axis_bram_74_tvalid(m_axis_bramio_74_tvalid),
        .m_axis_bram_74_tkeep(m_axis_bramio_74_tkeep),
        .m_axis_bram_74_tstrb(m_axis_bramio_74_tstrb),
        .m_axis_bram_74_tdata(m_axis_bramio_74_tdata),
        .m_axis_bram_74_tready(m_axis_bramio_74_tready),
        .m_axis_bram_75_tlast(m_axis_bramio_75_tlast),
        .m_axis_bram_75_tvalid(m_axis_bramio_75_tvalid),
        .m_axis_bram_75_tkeep(m_axis_bramio_75_tkeep),
        .m_axis_bram_75_tstrb(m_axis_bramio_75_tstrb),
        .m_axis_bram_75_tdata(m_axis_bramio_75_tdata),
        .m_axis_bram_75_tready(m_axis_bramio_75_tready),
        .m_axis_bram_76_tlast(m_axis_bramio_76_tlast),
        .m_axis_bram_76_tvalid(m_axis_bramio_76_tvalid),
        .m_axis_bram_76_tkeep(m_axis_bramio_76_tkeep),
        .m_axis_bram_76_tstrb(m_axis_bramio_76_tstrb),
        .m_axis_bram_76_tdata(m_axis_bramio_76_tdata),
        .m_axis_bram_76_tready(m_axis_bramio_76_tready),
        .m_axis_bram_77_tlast(m_axis_bramio_77_tlast),
        .m_axis_bram_77_tvalid(m_axis_bramio_77_tvalid),
        .m_axis_bram_77_tkeep(m_axis_bramio_77_tkeep),
        .m_axis_bram_77_tstrb(m_axis_bramio_77_tstrb),
        .m_axis_bram_77_tdata(m_axis_bramio_77_tdata),
        .m_axis_bram_77_tready(m_axis_bramio_77_tready),
        .m_axis_bram_78_tlast(m_axis_bramio_78_tlast),
        .m_axis_bram_78_tvalid(m_axis_bramio_78_tvalid),
        .m_axis_bram_78_tkeep(m_axis_bramio_78_tkeep),
        .m_axis_bram_78_tstrb(m_axis_bramio_78_tstrb),
        .m_axis_bram_78_tdata(m_axis_bramio_78_tdata),
        .m_axis_bram_78_tready(m_axis_bramio_78_tready),
        .m_axis_bram_79_tlast(m_axis_bramio_79_tlast),
        .m_axis_bram_79_tvalid(m_axis_bramio_79_tvalid),
        .m_axis_bram_79_tkeep(m_axis_bramio_79_tkeep),
        .m_axis_bram_79_tstrb(m_axis_bramio_79_tstrb),
        .m_axis_bram_79_tdata(m_axis_bramio_79_tdata),
        .m_axis_bram_79_tready(m_axis_bramio_79_tready),
        .m_axis_bram_80_tlast(m_axis_bramio_80_tlast),
        .m_axis_bram_80_tvalid(m_axis_bramio_80_tvalid),
        .m_axis_bram_80_tkeep(m_axis_bramio_80_tkeep),
        .m_axis_bram_80_tstrb(m_axis_bramio_80_tstrb),
        .m_axis_bram_80_tdata(m_axis_bramio_80_tdata),
        .m_axis_bram_80_tready(m_axis_bramio_80_tready),
        .m_axis_bram_81_tlast(m_axis_bramio_81_tlast),
        .m_axis_bram_81_tvalid(m_axis_bramio_81_tvalid),
        .m_axis_bram_81_tkeep(m_axis_bramio_81_tkeep),
        .m_axis_bram_81_tstrb(m_axis_bramio_81_tstrb),
        .m_axis_bram_81_tdata(m_axis_bramio_81_tdata),
        .m_axis_bram_81_tready(m_axis_bramio_81_tready),
        .m_axis_bram_82_tlast(m_axis_bramio_82_tlast),
        .m_axis_bram_82_tvalid(m_axis_bramio_82_tvalid),
        .m_axis_bram_82_tkeep(m_axis_bramio_82_tkeep),
        .m_axis_bram_82_tstrb(m_axis_bramio_82_tstrb),
        .m_axis_bram_82_tdata(m_axis_bramio_82_tdata),
        .m_axis_bram_82_tready(m_axis_bramio_82_tready),
        .m_axis_bram_83_tlast(m_axis_bramio_83_tlast),
        .m_axis_bram_83_tvalid(m_axis_bramio_83_tvalid),
        .m_axis_bram_83_tkeep(m_axis_bramio_83_tkeep),
        .m_axis_bram_83_tstrb(m_axis_bramio_83_tstrb),
        .m_axis_bram_83_tdata(m_axis_bramio_83_tdata),
        .m_axis_bram_83_tready(m_axis_bramio_83_tready),
        .m_axis_bram_84_tlast(m_axis_bramio_84_tlast),
        .m_axis_bram_84_tvalid(m_axis_bramio_84_tvalid),
        .m_axis_bram_84_tkeep(m_axis_bramio_84_tkeep),
        .m_axis_bram_84_tstrb(m_axis_bramio_84_tstrb),
        .m_axis_bram_84_tdata(m_axis_bramio_84_tdata),
        .m_axis_bram_84_tready(m_axis_bramio_84_tready),
        .m_axis_bram_85_tlast(m_axis_bramio_85_tlast),
        .m_axis_bram_85_tvalid(m_axis_bramio_85_tvalid),
        .m_axis_bram_85_tkeep(m_axis_bramio_85_tkeep),
        .m_axis_bram_85_tstrb(m_axis_bramio_85_tstrb),
        .m_axis_bram_85_tdata(m_axis_bramio_85_tdata),
        .m_axis_bram_85_tready(m_axis_bramio_85_tready),
        .m_axis_bram_86_tlast(m_axis_bramio_86_tlast),
        .m_axis_bram_86_tvalid(m_axis_bramio_86_tvalid),
        .m_axis_bram_86_tkeep(m_axis_bramio_86_tkeep),
        .m_axis_bram_86_tstrb(m_axis_bramio_86_tstrb),
        .m_axis_bram_86_tdata(m_axis_bramio_86_tdata),
        .m_axis_bram_86_tready(m_axis_bramio_86_tready),
        .m_axis_bram_87_tlast(m_axis_bramio_87_tlast),
        .m_axis_bram_87_tvalid(m_axis_bramio_87_tvalid),
        .m_axis_bram_87_tkeep(m_axis_bramio_87_tkeep),
        .m_axis_bram_87_tstrb(m_axis_bramio_87_tstrb),
        .m_axis_bram_87_tdata(m_axis_bramio_87_tdata),
        .m_axis_bram_87_tready(m_axis_bramio_87_tready),
        .m_axis_bram_88_tlast(m_axis_bramio_88_tlast),
        .m_axis_bram_88_tvalid(m_axis_bramio_88_tvalid),
        .m_axis_bram_88_tkeep(m_axis_bramio_88_tkeep),
        .m_axis_bram_88_tstrb(m_axis_bramio_88_tstrb),
        .m_axis_bram_88_tdata(m_axis_bramio_88_tdata),
        .m_axis_bram_88_tready(m_axis_bramio_88_tready),
        .m_axis_bram_89_tlast(m_axis_bramio_89_tlast),
        .m_axis_bram_89_tvalid(m_axis_bramio_89_tvalid),
        .m_axis_bram_89_tkeep(m_axis_bramio_89_tkeep),
        .m_axis_bram_89_tstrb(m_axis_bramio_89_tstrb),
        .m_axis_bram_89_tdata(m_axis_bramio_89_tdata),
        .m_axis_bram_89_tready(m_axis_bramio_89_tready),
        .m_axis_bram_90_tlast(m_axis_bramio_90_tlast),
        .m_axis_bram_90_tvalid(m_axis_bramio_90_tvalid),
        .m_axis_bram_90_tkeep(m_axis_bramio_90_tkeep),
        .m_axis_bram_90_tstrb(m_axis_bramio_90_tstrb),
        .m_axis_bram_90_tdata(m_axis_bramio_90_tdata),
        .m_axis_bram_90_tready(m_axis_bramio_90_tready),
        .m_axis_bram_91_tlast(m_axis_bramio_91_tlast),
        .m_axis_bram_91_tvalid(m_axis_bramio_91_tvalid),
        .m_axis_bram_91_tkeep(m_axis_bramio_91_tkeep),
        .m_axis_bram_91_tstrb(m_axis_bramio_91_tstrb),
        .m_axis_bram_91_tdata(m_axis_bramio_91_tdata),
        .m_axis_bram_91_tready(m_axis_bramio_91_tready),
        .m_axis_bram_92_tlast(m_axis_bramio_92_tlast),
        .m_axis_bram_92_tvalid(m_axis_bramio_92_tvalid),
        .m_axis_bram_92_tkeep(m_axis_bramio_92_tkeep),
        .m_axis_bram_92_tstrb(m_axis_bramio_92_tstrb),
        .m_axis_bram_92_tdata(m_axis_bramio_92_tdata),
        .m_axis_bram_92_tready(m_axis_bramio_92_tready),
        .m_axis_bram_93_tlast(m_axis_bramio_93_tlast),
        .m_axis_bram_93_tvalid(m_axis_bramio_93_tvalid),
        .m_axis_bram_93_tkeep(m_axis_bramio_93_tkeep),
        .m_axis_bram_93_tstrb(m_axis_bramio_93_tstrb),
        .m_axis_bram_93_tdata(m_axis_bramio_93_tdata),
        .m_axis_bram_93_tready(m_axis_bramio_93_tready),
        .m_axis_bram_94_tlast(m_axis_bramio_94_tlast),
        .m_axis_bram_94_tvalid(m_axis_bramio_94_tvalid),
        .m_axis_bram_94_tkeep(m_axis_bramio_94_tkeep),
        .m_axis_bram_94_tstrb(m_axis_bramio_94_tstrb),
        .m_axis_bram_94_tdata(m_axis_bramio_94_tdata),
        .m_axis_bram_94_tready(m_axis_bramio_94_tready),
        .m_axis_bram_95_tlast(m_axis_bramio_95_tlast),
        .m_axis_bram_95_tvalid(m_axis_bramio_95_tvalid),
        .m_axis_bram_95_tkeep(m_axis_bramio_95_tkeep),
        .m_axis_bram_95_tstrb(m_axis_bramio_95_tstrb),
        .m_axis_bram_95_tdata(m_axis_bramio_95_tdata),
        .m_axis_bram_95_tready(m_axis_bramio_95_tready),
        .m_axis_bram_96_tlast(m_axis_bramio_96_tlast),
        .m_axis_bram_96_tvalid(m_axis_bramio_96_tvalid),
        .m_axis_bram_96_tkeep(m_axis_bramio_96_tkeep),
        .m_axis_bram_96_tstrb(m_axis_bramio_96_tstrb),
        .m_axis_bram_96_tdata(m_axis_bramio_96_tdata),
        .m_axis_bram_96_tready(m_axis_bramio_96_tready),
        .m_axis_bram_97_tlast(m_axis_bramio_97_tlast),
        .m_axis_bram_97_tvalid(m_axis_bramio_97_tvalid),
        .m_axis_bram_97_tkeep(m_axis_bramio_97_tkeep),
        .m_axis_bram_97_tstrb(m_axis_bramio_97_tstrb),
        .m_axis_bram_97_tdata(m_axis_bramio_97_tdata),
        .m_axis_bram_97_tready(m_axis_bramio_97_tready),
        .m_axis_bram_98_tlast(m_axis_bramio_98_tlast),
        .m_axis_bram_98_tvalid(m_axis_bramio_98_tvalid),
        .m_axis_bram_98_tkeep(m_axis_bramio_98_tkeep),
        .m_axis_bram_98_tstrb(m_axis_bramio_98_tstrb),
        .m_axis_bram_98_tdata(m_axis_bramio_98_tdata),
        .m_axis_bram_98_tready(m_axis_bramio_98_tready),
        .m_axis_bram_99_tlast(m_axis_bramio_99_tlast),
        .m_axis_bram_99_tvalid(m_axis_bramio_99_tvalid),
        .m_axis_bram_99_tkeep(m_axis_bramio_99_tkeep),
        .m_axis_bram_99_tstrb(m_axis_bramio_99_tstrb),
        .m_axis_bram_99_tdata(m_axis_bramio_99_tdata),
        .m_axis_bram_99_tready(m_axis_bramio_99_tready),
        .m_axis_bram_100_tlast(m_axis_bramio_100_tlast),
        .m_axis_bram_100_tvalid(m_axis_bramio_100_tvalid),
        .m_axis_bram_100_tkeep(m_axis_bramio_100_tkeep),
        .m_axis_bram_100_tstrb(m_axis_bramio_100_tstrb),
        .m_axis_bram_100_tdata(m_axis_bramio_100_tdata),
        .m_axis_bram_100_tready(m_axis_bramio_100_tready),
        .m_axis_bram_101_tlast(m_axis_bramio_101_tlast),
        .m_axis_bram_101_tvalid(m_axis_bramio_101_tvalid),
        .m_axis_bram_101_tkeep(m_axis_bramio_101_tkeep),
        .m_axis_bram_101_tstrb(m_axis_bramio_101_tstrb),
        .m_axis_bram_101_tdata(m_axis_bramio_101_tdata),
        .m_axis_bram_101_tready(m_axis_bramio_101_tready),
        .m_axis_bram_102_tlast(m_axis_bramio_102_tlast),
        .m_axis_bram_102_tvalid(m_axis_bramio_102_tvalid),
        .m_axis_bram_102_tkeep(m_axis_bramio_102_tkeep),
        .m_axis_bram_102_tstrb(m_axis_bramio_102_tstrb),
        .m_axis_bram_102_tdata(m_axis_bramio_102_tdata),
        .m_axis_bram_102_tready(m_axis_bramio_102_tready),
        .m_axis_bram_103_tlast(m_axis_bramio_103_tlast),
        .m_axis_bram_103_tvalid(m_axis_bramio_103_tvalid),
        .m_axis_bram_103_tkeep(m_axis_bramio_103_tkeep),
        .m_axis_bram_103_tstrb(m_axis_bramio_103_tstrb),
        .m_axis_bram_103_tdata(m_axis_bramio_103_tdata),
        .m_axis_bram_103_tready(m_axis_bramio_103_tready),
        .m_axis_bram_104_tlast(m_axis_bramio_104_tlast),
        .m_axis_bram_104_tvalid(m_axis_bramio_104_tvalid),
        .m_axis_bram_104_tkeep(m_axis_bramio_104_tkeep),
        .m_axis_bram_104_tstrb(m_axis_bramio_104_tstrb),
        .m_axis_bram_104_tdata(m_axis_bramio_104_tdata),
        .m_axis_bram_104_tready(m_axis_bramio_104_tready),
        .m_axis_bram_105_tlast(m_axis_bramio_105_tlast),
        .m_axis_bram_105_tvalid(m_axis_bramio_105_tvalid),
        .m_axis_bram_105_tkeep(m_axis_bramio_105_tkeep),
        .m_axis_bram_105_tstrb(m_axis_bramio_105_tstrb),
        .m_axis_bram_105_tdata(m_axis_bramio_105_tdata),
        .m_axis_bram_105_tready(m_axis_bramio_105_tready),
        .m_axis_bram_106_tlast(m_axis_bramio_106_tlast),
        .m_axis_bram_106_tvalid(m_axis_bramio_106_tvalid),
        .m_axis_bram_106_tkeep(m_axis_bramio_106_tkeep),
        .m_axis_bram_106_tstrb(m_axis_bramio_106_tstrb),
        .m_axis_bram_106_tdata(m_axis_bramio_106_tdata),
        .m_axis_bram_106_tready(m_axis_bramio_106_tready),
        .m_axis_bram_107_tlast(m_axis_bramio_107_tlast),
        .m_axis_bram_107_tvalid(m_axis_bramio_107_tvalid),
        .m_axis_bram_107_tkeep(m_axis_bramio_107_tkeep),
        .m_axis_bram_107_tstrb(m_axis_bramio_107_tstrb),
        .m_axis_bram_107_tdata(m_axis_bramio_107_tdata),
        .m_axis_bram_107_tready(m_axis_bramio_107_tready),
        .m_axis_bram_108_tlast(m_axis_bramio_108_tlast),
        .m_axis_bram_108_tvalid(m_axis_bramio_108_tvalid),
        .m_axis_bram_108_tkeep(m_axis_bramio_108_tkeep),
        .m_axis_bram_108_tstrb(m_axis_bramio_108_tstrb),
        .m_axis_bram_108_tdata(m_axis_bramio_108_tdata),
        .m_axis_bram_108_tready(m_axis_bramio_108_tready),
        .m_axis_bram_109_tlast(m_axis_bramio_109_tlast),
        .m_axis_bram_109_tvalid(m_axis_bramio_109_tvalid),
        .m_axis_bram_109_tkeep(m_axis_bramio_109_tkeep),
        .m_axis_bram_109_tstrb(m_axis_bramio_109_tstrb),
        .m_axis_bram_109_tdata(m_axis_bramio_109_tdata),
        .m_axis_bram_109_tready(m_axis_bramio_109_tready),
        .m_axis_bram_110_tlast(m_axis_bramio_110_tlast),
        .m_axis_bram_110_tvalid(m_axis_bramio_110_tvalid),
        .m_axis_bram_110_tkeep(m_axis_bramio_110_tkeep),
        .m_axis_bram_110_tstrb(m_axis_bramio_110_tstrb),
        .m_axis_bram_110_tdata(m_axis_bramio_110_tdata),
        .m_axis_bram_110_tready(m_axis_bramio_110_tready),
        .m_axis_bram_111_tlast(m_axis_bramio_111_tlast),
        .m_axis_bram_111_tvalid(m_axis_bramio_111_tvalid),
        .m_axis_bram_111_tkeep(m_axis_bramio_111_tkeep),
        .m_axis_bram_111_tstrb(m_axis_bramio_111_tstrb),
        .m_axis_bram_111_tdata(m_axis_bramio_111_tdata),
        .m_axis_bram_111_tready(m_axis_bramio_111_tready),
        .m_axis_bram_112_tlast(m_axis_bramio_112_tlast),
        .m_axis_bram_112_tvalid(m_axis_bramio_112_tvalid),
        .m_axis_bram_112_tkeep(m_axis_bramio_112_tkeep),
        .m_axis_bram_112_tstrb(m_axis_bramio_112_tstrb),
        .m_axis_bram_112_tdata(m_axis_bramio_112_tdata),
        .m_axis_bram_112_tready(m_axis_bramio_112_tready),
        .m_axis_bram_113_tlast(m_axis_bramio_113_tlast),
        .m_axis_bram_113_tvalid(m_axis_bramio_113_tvalid),
        .m_axis_bram_113_tkeep(m_axis_bramio_113_tkeep),
        .m_axis_bram_113_tstrb(m_axis_bramio_113_tstrb),
        .m_axis_bram_113_tdata(m_axis_bramio_113_tdata),
        .m_axis_bram_113_tready(m_axis_bramio_113_tready),
        .m_axis_bram_114_tlast(m_axis_bramio_114_tlast),
        .m_axis_bram_114_tvalid(m_axis_bramio_114_tvalid),
        .m_axis_bram_114_tkeep(m_axis_bramio_114_tkeep),
        .m_axis_bram_114_tstrb(m_axis_bramio_114_tstrb),
        .m_axis_bram_114_tdata(m_axis_bramio_114_tdata),
        .m_axis_bram_114_tready(m_axis_bramio_114_tready),
        .m_axis_bram_115_tlast(m_axis_bramio_115_tlast),
        .m_axis_bram_115_tvalid(m_axis_bramio_115_tvalid),
        .m_axis_bram_115_tkeep(m_axis_bramio_115_tkeep),
        .m_axis_bram_115_tstrb(m_axis_bramio_115_tstrb),
        .m_axis_bram_115_tdata(m_axis_bramio_115_tdata),
        .m_axis_bram_115_tready(m_axis_bramio_115_tready),
        .m_axis_bram_116_tlast(m_axis_bramio_116_tlast),
        .m_axis_bram_116_tvalid(m_axis_bramio_116_tvalid),
        .m_axis_bram_116_tkeep(m_axis_bramio_116_tkeep),
        .m_axis_bram_116_tstrb(m_axis_bramio_116_tstrb),
        .m_axis_bram_116_tdata(m_axis_bramio_116_tdata),
        .m_axis_bram_116_tready(m_axis_bramio_116_tready),
        .m_axis_bram_117_tlast(m_axis_bramio_117_tlast),
        .m_axis_bram_117_tvalid(m_axis_bramio_117_tvalid),
        .m_axis_bram_117_tkeep(m_axis_bramio_117_tkeep),
        .m_axis_bram_117_tstrb(m_axis_bramio_117_tstrb),
        .m_axis_bram_117_tdata(m_axis_bramio_117_tdata),
        .m_axis_bram_117_tready(m_axis_bramio_117_tready),
        .m_axis_bram_118_tlast(m_axis_bramio_118_tlast),
        .m_axis_bram_118_tvalid(m_axis_bramio_118_tvalid),
        .m_axis_bram_118_tkeep(m_axis_bramio_118_tkeep),
        .m_axis_bram_118_tstrb(m_axis_bramio_118_tstrb),
        .m_axis_bram_118_tdata(m_axis_bramio_118_tdata),
        .m_axis_bram_118_tready(m_axis_bramio_118_tready),
        .m_axis_bram_119_tlast(m_axis_bramio_119_tlast),
        .m_axis_bram_119_tvalid(m_axis_bramio_119_tvalid),
        .m_axis_bram_119_tkeep(m_axis_bramio_119_tkeep),
        .m_axis_bram_119_tstrb(m_axis_bramio_119_tstrb),
        .m_axis_bram_119_tdata(m_axis_bramio_119_tdata),
        .m_axis_bram_119_tready(m_axis_bramio_119_tready),
        .m_axis_bram_120_tlast(m_axis_bramio_120_tlast),
        .m_axis_bram_120_tvalid(m_axis_bramio_120_tvalid),
        .m_axis_bram_120_tkeep(m_axis_bramio_120_tkeep),
        .m_axis_bram_120_tstrb(m_axis_bramio_120_tstrb),
        .m_axis_bram_120_tdata(m_axis_bramio_120_tdata),
        .m_axis_bram_120_tready(m_axis_bramio_120_tready),
        .m_axis_bram_121_tlast(m_axis_bramio_121_tlast),
        .m_axis_bram_121_tvalid(m_axis_bramio_121_tvalid),
        .m_axis_bram_121_tkeep(m_axis_bramio_121_tkeep),
        .m_axis_bram_121_tstrb(m_axis_bramio_121_tstrb),
        .m_axis_bram_121_tdata(m_axis_bramio_121_tdata),
        .m_axis_bram_121_tready(m_axis_bramio_121_tready),
        .m_axis_bram_122_tlast(m_axis_bramio_122_tlast),
        .m_axis_bram_122_tvalid(m_axis_bramio_122_tvalid),
        .m_axis_bram_122_tkeep(m_axis_bramio_122_tkeep),
        .m_axis_bram_122_tstrb(m_axis_bramio_122_tstrb),
        .m_axis_bram_122_tdata(m_axis_bramio_122_tdata),
        .m_axis_bram_122_tready(m_axis_bramio_122_tready),
        .m_axis_bram_123_tlast(m_axis_bramio_123_tlast),
        .m_axis_bram_123_tvalid(m_axis_bramio_123_tvalid),
        .m_axis_bram_123_tkeep(m_axis_bramio_123_tkeep),
        .m_axis_bram_123_tstrb(m_axis_bramio_123_tstrb),
        .m_axis_bram_123_tdata(m_axis_bramio_123_tdata),
        .m_axis_bram_123_tready(m_axis_bramio_123_tready),
        .m_axis_bram_124_tlast(m_axis_bramio_124_tlast),
        .m_axis_bram_124_tvalid(m_axis_bramio_124_tvalid),
        .m_axis_bram_124_tkeep(m_axis_bramio_124_tkeep),
        .m_axis_bram_124_tstrb(m_axis_bramio_124_tstrb),
        .m_axis_bram_124_tdata(m_axis_bramio_124_tdata),
        .m_axis_bram_124_tready(m_axis_bramio_124_tready),
        .m_axis_bram_125_tlast(m_axis_bramio_125_tlast),
        .m_axis_bram_125_tvalid(m_axis_bramio_125_tvalid),
        .m_axis_bram_125_tkeep(m_axis_bramio_125_tkeep),
        .m_axis_bram_125_tstrb(m_axis_bramio_125_tstrb),
        .m_axis_bram_125_tdata(m_axis_bramio_125_tdata),
        .m_axis_bram_125_tready(m_axis_bramio_125_tready),
        .m_axis_bram_126_tlast(m_axis_bramio_126_tlast),
        .m_axis_bram_126_tvalid(m_axis_bramio_126_tvalid),
        .m_axis_bram_126_tkeep(m_axis_bramio_126_tkeep),
        .m_axis_bram_126_tstrb(m_axis_bramio_126_tstrb),
        .m_axis_bram_126_tdata(m_axis_bramio_126_tdata),
        .m_axis_bram_126_tready(m_axis_bramio_126_tready),
        .m_axis_bram_127_tlast(m_axis_bramio_127_tlast),
        .m_axis_bram_127_tvalid(m_axis_bramio_127_tvalid),
        .m_axis_bram_127_tkeep(m_axis_bramio_127_tkeep),
        .m_axis_bram_127_tstrb(m_axis_bramio_127_tstrb),
        .m_axis_bram_127_tdata(m_axis_bramio_127_tdata),
        .m_axis_bram_127_tready(m_axis_bramio_127_tready)
    );
    
    out_bram_args #(
        .C_QUEUE_DEPTH(C_QUEUE_DEPTH),
        .C_NUM_OUTPUT_BRAMs(C_NUM_OUTPUT_BRAMs),
        .C_OUTPUT_BRAM_0_WIDTH(C_OUTPUT_BRAM_0_WIDTH),
        .C_OUTPUT_BRAM_1_WIDTH(C_OUTPUT_BRAM_1_WIDTH),
        .C_OUTPUT_BRAM_2_WIDTH(C_OUTPUT_BRAM_2_WIDTH),
        .C_OUTPUT_BRAM_3_WIDTH(C_OUTPUT_BRAM_3_WIDTH),
        .C_OUTPUT_BRAM_4_WIDTH(C_OUTPUT_BRAM_4_WIDTH),
        .C_OUTPUT_BRAM_5_WIDTH(C_OUTPUT_BRAM_5_WIDTH),
        .C_OUTPUT_BRAM_6_WIDTH(C_OUTPUT_BRAM_6_WIDTH),
        .C_OUTPUT_BRAM_7_WIDTH(C_OUTPUT_BRAM_7_WIDTH),
        .C_OUTPUT_BRAM_8_WIDTH(C_OUTPUT_BRAM_8_WIDTH),
        .C_OUTPUT_BRAM_9_WIDTH(C_OUTPUT_BRAM_9_WIDTH),
        .C_OUTPUT_BRAM_10_WIDTH(C_OUTPUT_BRAM_10_WIDTH),
        .C_OUTPUT_BRAM_11_WIDTH(C_OUTPUT_BRAM_11_WIDTH),
        .C_OUTPUT_BRAM_12_WIDTH(C_OUTPUT_BRAM_12_WIDTH),
        .C_OUTPUT_BRAM_13_WIDTH(C_OUTPUT_BRAM_13_WIDTH),
        .C_OUTPUT_BRAM_14_WIDTH(C_OUTPUT_BRAM_14_WIDTH),
        .C_OUTPUT_BRAM_15_WIDTH(C_OUTPUT_BRAM_15_WIDTH),
        .C_OUTPUT_BRAM_16_WIDTH(C_OUTPUT_BRAM_16_WIDTH),
        .C_OUTPUT_BRAM_17_WIDTH(C_OUTPUT_BRAM_17_WIDTH),
        .C_OUTPUT_BRAM_18_WIDTH(C_OUTPUT_BRAM_18_WIDTH),
        .C_OUTPUT_BRAM_19_WIDTH(C_OUTPUT_BRAM_19_WIDTH),
        .C_OUTPUT_BRAM_20_WIDTH(C_OUTPUT_BRAM_20_WIDTH),
        .C_OUTPUT_BRAM_21_WIDTH(C_OUTPUT_BRAM_21_WIDTH),
        .C_OUTPUT_BRAM_22_WIDTH(C_OUTPUT_BRAM_22_WIDTH),
        .C_OUTPUT_BRAM_23_WIDTH(C_OUTPUT_BRAM_23_WIDTH),
        .C_OUTPUT_BRAM_24_WIDTH(C_OUTPUT_BRAM_24_WIDTH),
        .C_OUTPUT_BRAM_25_WIDTH(C_OUTPUT_BRAM_25_WIDTH),
        .C_OUTPUT_BRAM_26_WIDTH(C_OUTPUT_BRAM_26_WIDTH),
        .C_OUTPUT_BRAM_27_WIDTH(C_OUTPUT_BRAM_27_WIDTH),
        .C_OUTPUT_BRAM_28_WIDTH(C_OUTPUT_BRAM_28_WIDTH),
        .C_OUTPUT_BRAM_29_WIDTH(C_OUTPUT_BRAM_29_WIDTH),
        .C_OUTPUT_BRAM_30_WIDTH(C_OUTPUT_BRAM_30_WIDTH),
        .C_OUTPUT_BRAM_31_WIDTH(C_OUTPUT_BRAM_31_WIDTH),
        .C_OUTPUT_BRAM_32_WIDTH(C_OUTPUT_BRAM_32_WIDTH),
        .C_OUTPUT_BRAM_33_WIDTH(C_OUTPUT_BRAM_33_WIDTH),
        .C_OUTPUT_BRAM_34_WIDTH(C_OUTPUT_BRAM_34_WIDTH),
        .C_OUTPUT_BRAM_35_WIDTH(C_OUTPUT_BRAM_35_WIDTH),
        .C_OUTPUT_BRAM_36_WIDTH(C_OUTPUT_BRAM_36_WIDTH),
        .C_OUTPUT_BRAM_37_WIDTH(C_OUTPUT_BRAM_37_WIDTH),
        .C_OUTPUT_BRAM_38_WIDTH(C_OUTPUT_BRAM_38_WIDTH),
        .C_OUTPUT_BRAM_39_WIDTH(C_OUTPUT_BRAM_39_WIDTH),
        .C_OUTPUT_BRAM_40_WIDTH(C_OUTPUT_BRAM_40_WIDTH),
        .C_OUTPUT_BRAM_41_WIDTH(C_OUTPUT_BRAM_41_WIDTH),
        .C_OUTPUT_BRAM_42_WIDTH(C_OUTPUT_BRAM_42_WIDTH),
        .C_OUTPUT_BRAM_43_WIDTH(C_OUTPUT_BRAM_43_WIDTH),
        .C_OUTPUT_BRAM_44_WIDTH(C_OUTPUT_BRAM_44_WIDTH),
        .C_OUTPUT_BRAM_45_WIDTH(C_OUTPUT_BRAM_45_WIDTH),
        .C_OUTPUT_BRAM_46_WIDTH(C_OUTPUT_BRAM_46_WIDTH),
        .C_OUTPUT_BRAM_47_WIDTH(C_OUTPUT_BRAM_47_WIDTH),
        .C_OUTPUT_BRAM_48_WIDTH(C_OUTPUT_BRAM_48_WIDTH),
        .C_OUTPUT_BRAM_49_WIDTH(C_OUTPUT_BRAM_49_WIDTH),
        .C_OUTPUT_BRAM_50_WIDTH(C_OUTPUT_BRAM_50_WIDTH),
        .C_OUTPUT_BRAM_51_WIDTH(C_OUTPUT_BRAM_51_WIDTH),
        .C_OUTPUT_BRAM_52_WIDTH(C_OUTPUT_BRAM_52_WIDTH),
        .C_OUTPUT_BRAM_53_WIDTH(C_OUTPUT_BRAM_53_WIDTH),
        .C_OUTPUT_BRAM_54_WIDTH(C_OUTPUT_BRAM_54_WIDTH),
        .C_OUTPUT_BRAM_55_WIDTH(C_OUTPUT_BRAM_55_WIDTH),
        .C_OUTPUT_BRAM_56_WIDTH(C_OUTPUT_BRAM_56_WIDTH),
        .C_OUTPUT_BRAM_57_WIDTH(C_OUTPUT_BRAM_57_WIDTH),
        .C_OUTPUT_BRAM_58_WIDTH(C_OUTPUT_BRAM_58_WIDTH),
        .C_OUTPUT_BRAM_59_WIDTH(C_OUTPUT_BRAM_59_WIDTH),
        .C_OUTPUT_BRAM_60_WIDTH(C_OUTPUT_BRAM_60_WIDTH),
        .C_OUTPUT_BRAM_61_WIDTH(C_OUTPUT_BRAM_61_WIDTH),
        .C_OUTPUT_BRAM_62_WIDTH(C_OUTPUT_BRAM_62_WIDTH),
        .C_OUTPUT_BRAM_63_WIDTH(C_OUTPUT_BRAM_63_WIDTH),
        .C_OUTPUT_BRAM_64_WIDTH(C_OUTPUT_BRAM_64_WIDTH),
        .C_OUTPUT_BRAM_65_WIDTH(C_OUTPUT_BRAM_65_WIDTH),
        .C_OUTPUT_BRAM_66_WIDTH(C_OUTPUT_BRAM_66_WIDTH),
        .C_OUTPUT_BRAM_67_WIDTH(C_OUTPUT_BRAM_67_WIDTH),
        .C_OUTPUT_BRAM_68_WIDTH(C_OUTPUT_BRAM_68_WIDTH),
        .C_OUTPUT_BRAM_69_WIDTH(C_OUTPUT_BRAM_69_WIDTH),
        .C_OUTPUT_BRAM_70_WIDTH(C_OUTPUT_BRAM_70_WIDTH),
        .C_OUTPUT_BRAM_71_WIDTH(C_OUTPUT_BRAM_71_WIDTH),
        .C_OUTPUT_BRAM_72_WIDTH(C_OUTPUT_BRAM_72_WIDTH),
        .C_OUTPUT_BRAM_73_WIDTH(C_OUTPUT_BRAM_73_WIDTH),
        .C_OUTPUT_BRAM_74_WIDTH(C_OUTPUT_BRAM_74_WIDTH),
        .C_OUTPUT_BRAM_75_WIDTH(C_OUTPUT_BRAM_75_WIDTH),
        .C_OUTPUT_BRAM_76_WIDTH(C_OUTPUT_BRAM_76_WIDTH),
        .C_OUTPUT_BRAM_77_WIDTH(C_OUTPUT_BRAM_77_WIDTH),
        .C_OUTPUT_BRAM_78_WIDTH(C_OUTPUT_BRAM_78_WIDTH),
        .C_OUTPUT_BRAM_79_WIDTH(C_OUTPUT_BRAM_79_WIDTH),
        .C_OUTPUT_BRAM_80_WIDTH(C_OUTPUT_BRAM_80_WIDTH),
        .C_OUTPUT_BRAM_81_WIDTH(C_OUTPUT_BRAM_81_WIDTH),
        .C_OUTPUT_BRAM_82_WIDTH(C_OUTPUT_BRAM_82_WIDTH),
        .C_OUTPUT_BRAM_83_WIDTH(C_OUTPUT_BRAM_83_WIDTH),
        .C_OUTPUT_BRAM_84_WIDTH(C_OUTPUT_BRAM_84_WIDTH),
        .C_OUTPUT_BRAM_85_WIDTH(C_OUTPUT_BRAM_85_WIDTH),
        .C_OUTPUT_BRAM_86_WIDTH(C_OUTPUT_BRAM_86_WIDTH),
        .C_OUTPUT_BRAM_87_WIDTH(C_OUTPUT_BRAM_87_WIDTH),
        .C_OUTPUT_BRAM_88_WIDTH(C_OUTPUT_BRAM_88_WIDTH),
        .C_OUTPUT_BRAM_89_WIDTH(C_OUTPUT_BRAM_89_WIDTH),
        .C_OUTPUT_BRAM_90_WIDTH(C_OUTPUT_BRAM_90_WIDTH),
        .C_OUTPUT_BRAM_91_WIDTH(C_OUTPUT_BRAM_91_WIDTH),
        .C_OUTPUT_BRAM_92_WIDTH(C_OUTPUT_BRAM_92_WIDTH),
        .C_OUTPUT_BRAM_93_WIDTH(C_OUTPUT_BRAM_93_WIDTH),
        .C_OUTPUT_BRAM_94_WIDTH(C_OUTPUT_BRAM_94_WIDTH),
        .C_OUTPUT_BRAM_95_WIDTH(C_OUTPUT_BRAM_95_WIDTH),
        .C_OUTPUT_BRAM_96_WIDTH(C_OUTPUT_BRAM_96_WIDTH),
        .C_OUTPUT_BRAM_97_WIDTH(C_OUTPUT_BRAM_97_WIDTH),
        .C_OUTPUT_BRAM_98_WIDTH(C_OUTPUT_BRAM_98_WIDTH),
        .C_OUTPUT_BRAM_99_WIDTH(C_OUTPUT_BRAM_99_WIDTH),
        .C_OUTPUT_BRAM_100_WIDTH(C_OUTPUT_BRAM_100_WIDTH),
        .C_OUTPUT_BRAM_101_WIDTH(C_OUTPUT_BRAM_101_WIDTH),
        .C_OUTPUT_BRAM_102_WIDTH(C_OUTPUT_BRAM_102_WIDTH),
        .C_OUTPUT_BRAM_103_WIDTH(C_OUTPUT_BRAM_103_WIDTH),
        .C_OUTPUT_BRAM_104_WIDTH(C_OUTPUT_BRAM_104_WIDTH),
        .C_OUTPUT_BRAM_105_WIDTH(C_OUTPUT_BRAM_105_WIDTH),
        .C_OUTPUT_BRAM_106_WIDTH(C_OUTPUT_BRAM_106_WIDTH),
        .C_OUTPUT_BRAM_107_WIDTH(C_OUTPUT_BRAM_107_WIDTH),
        .C_OUTPUT_BRAM_108_WIDTH(C_OUTPUT_BRAM_108_WIDTH),
        .C_OUTPUT_BRAM_109_WIDTH(C_OUTPUT_BRAM_109_WIDTH),
        .C_OUTPUT_BRAM_110_WIDTH(C_OUTPUT_BRAM_110_WIDTH),
        .C_OUTPUT_BRAM_111_WIDTH(C_OUTPUT_BRAM_111_WIDTH),
        .C_OUTPUT_BRAM_112_WIDTH(C_OUTPUT_BRAM_112_WIDTH),
        .C_OUTPUT_BRAM_113_WIDTH(C_OUTPUT_BRAM_113_WIDTH),
        .C_OUTPUT_BRAM_114_WIDTH(C_OUTPUT_BRAM_114_WIDTH),
        .C_OUTPUT_BRAM_115_WIDTH(C_OUTPUT_BRAM_115_WIDTH),
        .C_OUTPUT_BRAM_116_WIDTH(C_OUTPUT_BRAM_116_WIDTH),
        .C_OUTPUT_BRAM_117_WIDTH(C_OUTPUT_BRAM_117_WIDTH),
        .C_OUTPUT_BRAM_118_WIDTH(C_OUTPUT_BRAM_118_WIDTH),
        .C_OUTPUT_BRAM_119_WIDTH(C_OUTPUT_BRAM_119_WIDTH),
        .C_OUTPUT_BRAM_120_WIDTH(C_OUTPUT_BRAM_120_WIDTH),
        .C_OUTPUT_BRAM_121_WIDTH(C_OUTPUT_BRAM_121_WIDTH),
        .C_OUTPUT_BRAM_122_WIDTH(C_OUTPUT_BRAM_122_WIDTH),
        .C_OUTPUT_BRAM_123_WIDTH(C_OUTPUT_BRAM_123_WIDTH),
        .C_OUTPUT_BRAM_124_WIDTH(C_OUTPUT_BRAM_124_WIDTH),
        .C_OUTPUT_BRAM_125_WIDTH(C_OUTPUT_BRAM_125_WIDTH),
        .C_OUTPUT_BRAM_126_WIDTH(C_OUTPUT_BRAM_126_WIDTH),
        .C_OUTPUT_BRAM_127_WIDTH(C_OUTPUT_BRAM_127_WIDTH),
        .C_OUTPUT_BRAM_0_DEPTH(C_OUTPUT_BRAM_0_DEPTH),
        .C_OUTPUT_BRAM_1_DEPTH(C_OUTPUT_BRAM_1_DEPTH),
        .C_OUTPUT_BRAM_2_DEPTH(C_OUTPUT_BRAM_2_DEPTH),
        .C_OUTPUT_BRAM_3_DEPTH(C_OUTPUT_BRAM_3_DEPTH),
        .C_OUTPUT_BRAM_4_DEPTH(C_OUTPUT_BRAM_4_DEPTH),
        .C_OUTPUT_BRAM_5_DEPTH(C_OUTPUT_BRAM_5_DEPTH),
        .C_OUTPUT_BRAM_6_DEPTH(C_OUTPUT_BRAM_6_DEPTH),
        .C_OUTPUT_BRAM_7_DEPTH(C_OUTPUT_BRAM_7_DEPTH),
        .C_OUTPUT_BRAM_8_DEPTH(C_OUTPUT_BRAM_8_DEPTH),
        .C_OUTPUT_BRAM_9_DEPTH(C_OUTPUT_BRAM_9_DEPTH),
        .C_OUTPUT_BRAM_10_DEPTH(C_OUTPUT_BRAM_10_DEPTH),
        .C_OUTPUT_BRAM_11_DEPTH(C_OUTPUT_BRAM_11_DEPTH),
        .C_OUTPUT_BRAM_12_DEPTH(C_OUTPUT_BRAM_12_DEPTH),
        .C_OUTPUT_BRAM_13_DEPTH(C_OUTPUT_BRAM_13_DEPTH),
        .C_OUTPUT_BRAM_14_DEPTH(C_OUTPUT_BRAM_14_DEPTH),
        .C_OUTPUT_BRAM_15_DEPTH(C_OUTPUT_BRAM_15_DEPTH),
        .C_OUTPUT_BRAM_16_DEPTH(C_OUTPUT_BRAM_16_DEPTH),
        .C_OUTPUT_BRAM_17_DEPTH(C_OUTPUT_BRAM_17_DEPTH),
        .C_OUTPUT_BRAM_18_DEPTH(C_OUTPUT_BRAM_18_DEPTH),
        .C_OUTPUT_BRAM_19_DEPTH(C_OUTPUT_BRAM_19_DEPTH),
        .C_OUTPUT_BRAM_20_DEPTH(C_OUTPUT_BRAM_20_DEPTH),
        .C_OUTPUT_BRAM_21_DEPTH(C_OUTPUT_BRAM_21_DEPTH),
        .C_OUTPUT_BRAM_22_DEPTH(C_OUTPUT_BRAM_22_DEPTH),
        .C_OUTPUT_BRAM_23_DEPTH(C_OUTPUT_BRAM_23_DEPTH),
        .C_OUTPUT_BRAM_24_DEPTH(C_OUTPUT_BRAM_24_DEPTH),
        .C_OUTPUT_BRAM_25_DEPTH(C_OUTPUT_BRAM_25_DEPTH),
        .C_OUTPUT_BRAM_26_DEPTH(C_OUTPUT_BRAM_26_DEPTH),
        .C_OUTPUT_BRAM_27_DEPTH(C_OUTPUT_BRAM_27_DEPTH),
        .C_OUTPUT_BRAM_28_DEPTH(C_OUTPUT_BRAM_28_DEPTH),
        .C_OUTPUT_BRAM_29_DEPTH(C_OUTPUT_BRAM_29_DEPTH),
        .C_OUTPUT_BRAM_30_DEPTH(C_OUTPUT_BRAM_30_DEPTH),
        .C_OUTPUT_BRAM_31_DEPTH(C_OUTPUT_BRAM_31_DEPTH),
        .C_OUTPUT_BRAM_32_DEPTH(C_OUTPUT_BRAM_32_DEPTH),
        .C_OUTPUT_BRAM_33_DEPTH(C_OUTPUT_BRAM_33_DEPTH),
        .C_OUTPUT_BRAM_34_DEPTH(C_OUTPUT_BRAM_34_DEPTH),
        .C_OUTPUT_BRAM_35_DEPTH(C_OUTPUT_BRAM_35_DEPTH),
        .C_OUTPUT_BRAM_36_DEPTH(C_OUTPUT_BRAM_36_DEPTH),
        .C_OUTPUT_BRAM_37_DEPTH(C_OUTPUT_BRAM_37_DEPTH),
        .C_OUTPUT_BRAM_38_DEPTH(C_OUTPUT_BRAM_38_DEPTH),
        .C_OUTPUT_BRAM_39_DEPTH(C_OUTPUT_BRAM_39_DEPTH),
        .C_OUTPUT_BRAM_40_DEPTH(C_OUTPUT_BRAM_40_DEPTH),
        .C_OUTPUT_BRAM_41_DEPTH(C_OUTPUT_BRAM_41_DEPTH),
        .C_OUTPUT_BRAM_42_DEPTH(C_OUTPUT_BRAM_42_DEPTH),
        .C_OUTPUT_BRAM_43_DEPTH(C_OUTPUT_BRAM_43_DEPTH),
        .C_OUTPUT_BRAM_44_DEPTH(C_OUTPUT_BRAM_44_DEPTH),
        .C_OUTPUT_BRAM_45_DEPTH(C_OUTPUT_BRAM_45_DEPTH),
        .C_OUTPUT_BRAM_46_DEPTH(C_OUTPUT_BRAM_46_DEPTH),
        .C_OUTPUT_BRAM_47_DEPTH(C_OUTPUT_BRAM_47_DEPTH),
        .C_OUTPUT_BRAM_48_DEPTH(C_OUTPUT_BRAM_48_DEPTH),
        .C_OUTPUT_BRAM_49_DEPTH(C_OUTPUT_BRAM_49_DEPTH),
        .C_OUTPUT_BRAM_50_DEPTH(C_OUTPUT_BRAM_50_DEPTH),
        .C_OUTPUT_BRAM_51_DEPTH(C_OUTPUT_BRAM_51_DEPTH),
        .C_OUTPUT_BRAM_52_DEPTH(C_OUTPUT_BRAM_52_DEPTH),
        .C_OUTPUT_BRAM_53_DEPTH(C_OUTPUT_BRAM_53_DEPTH),
        .C_OUTPUT_BRAM_54_DEPTH(C_OUTPUT_BRAM_54_DEPTH),
        .C_OUTPUT_BRAM_55_DEPTH(C_OUTPUT_BRAM_55_DEPTH),
        .C_OUTPUT_BRAM_56_DEPTH(C_OUTPUT_BRAM_56_DEPTH),
        .C_OUTPUT_BRAM_57_DEPTH(C_OUTPUT_BRAM_57_DEPTH),
        .C_OUTPUT_BRAM_58_DEPTH(C_OUTPUT_BRAM_58_DEPTH),
        .C_OUTPUT_BRAM_59_DEPTH(C_OUTPUT_BRAM_59_DEPTH),
        .C_OUTPUT_BRAM_60_DEPTH(C_OUTPUT_BRAM_60_DEPTH),
        .C_OUTPUT_BRAM_61_DEPTH(C_OUTPUT_BRAM_61_DEPTH),
        .C_OUTPUT_BRAM_62_DEPTH(C_OUTPUT_BRAM_62_DEPTH),
        .C_OUTPUT_BRAM_63_DEPTH(C_OUTPUT_BRAM_63_DEPTH),
        .C_OUTPUT_BRAM_64_DEPTH(C_OUTPUT_BRAM_64_DEPTH),
        .C_OUTPUT_BRAM_65_DEPTH(C_OUTPUT_BRAM_65_DEPTH),
        .C_OUTPUT_BRAM_66_DEPTH(C_OUTPUT_BRAM_66_DEPTH),
        .C_OUTPUT_BRAM_67_DEPTH(C_OUTPUT_BRAM_67_DEPTH),
        .C_OUTPUT_BRAM_68_DEPTH(C_OUTPUT_BRAM_68_DEPTH),
        .C_OUTPUT_BRAM_69_DEPTH(C_OUTPUT_BRAM_69_DEPTH),
        .C_OUTPUT_BRAM_70_DEPTH(C_OUTPUT_BRAM_70_DEPTH),
        .C_OUTPUT_BRAM_71_DEPTH(C_OUTPUT_BRAM_71_DEPTH),
        .C_OUTPUT_BRAM_72_DEPTH(C_OUTPUT_BRAM_72_DEPTH),
        .C_OUTPUT_BRAM_73_DEPTH(C_OUTPUT_BRAM_73_DEPTH),
        .C_OUTPUT_BRAM_74_DEPTH(C_OUTPUT_BRAM_74_DEPTH),
        .C_OUTPUT_BRAM_75_DEPTH(C_OUTPUT_BRAM_75_DEPTH),
        .C_OUTPUT_BRAM_76_DEPTH(C_OUTPUT_BRAM_76_DEPTH),
        .C_OUTPUT_BRAM_77_DEPTH(C_OUTPUT_BRAM_77_DEPTH),
        .C_OUTPUT_BRAM_78_DEPTH(C_OUTPUT_BRAM_78_DEPTH),
        .C_OUTPUT_BRAM_79_DEPTH(C_OUTPUT_BRAM_79_DEPTH),
        .C_OUTPUT_BRAM_80_DEPTH(C_OUTPUT_BRAM_80_DEPTH),
        .C_OUTPUT_BRAM_81_DEPTH(C_OUTPUT_BRAM_81_DEPTH),
        .C_OUTPUT_BRAM_82_DEPTH(C_OUTPUT_BRAM_82_DEPTH),
        .C_OUTPUT_BRAM_83_DEPTH(C_OUTPUT_BRAM_83_DEPTH),
        .C_OUTPUT_BRAM_84_DEPTH(C_OUTPUT_BRAM_84_DEPTH),
        .C_OUTPUT_BRAM_85_DEPTH(C_OUTPUT_BRAM_85_DEPTH),
        .C_OUTPUT_BRAM_86_DEPTH(C_OUTPUT_BRAM_86_DEPTH),
        .C_OUTPUT_BRAM_87_DEPTH(C_OUTPUT_BRAM_87_DEPTH),
        .C_OUTPUT_BRAM_88_DEPTH(C_OUTPUT_BRAM_88_DEPTH),
        .C_OUTPUT_BRAM_89_DEPTH(C_OUTPUT_BRAM_89_DEPTH),
        .C_OUTPUT_BRAM_90_DEPTH(C_OUTPUT_BRAM_90_DEPTH),
        .C_OUTPUT_BRAM_91_DEPTH(C_OUTPUT_BRAM_91_DEPTH),
        .C_OUTPUT_BRAM_92_DEPTH(C_OUTPUT_BRAM_92_DEPTH),
        .C_OUTPUT_BRAM_93_DEPTH(C_OUTPUT_BRAM_93_DEPTH),
        .C_OUTPUT_BRAM_94_DEPTH(C_OUTPUT_BRAM_94_DEPTH),
        .C_OUTPUT_BRAM_95_DEPTH(C_OUTPUT_BRAM_95_DEPTH),
        .C_OUTPUT_BRAM_96_DEPTH(C_OUTPUT_BRAM_96_DEPTH),
        .C_OUTPUT_BRAM_97_DEPTH(C_OUTPUT_BRAM_97_DEPTH),
        .C_OUTPUT_BRAM_98_DEPTH(C_OUTPUT_BRAM_98_DEPTH),
        .C_OUTPUT_BRAM_99_DEPTH(C_OUTPUT_BRAM_99_DEPTH),
        .C_OUTPUT_BRAM_100_DEPTH(C_OUTPUT_BRAM_100_DEPTH),
        .C_OUTPUT_BRAM_101_DEPTH(C_OUTPUT_BRAM_101_DEPTH),
        .C_OUTPUT_BRAM_102_DEPTH(C_OUTPUT_BRAM_102_DEPTH),
        .C_OUTPUT_BRAM_103_DEPTH(C_OUTPUT_BRAM_103_DEPTH),
        .C_OUTPUT_BRAM_104_DEPTH(C_OUTPUT_BRAM_104_DEPTH),
        .C_OUTPUT_BRAM_105_DEPTH(C_OUTPUT_BRAM_105_DEPTH),
        .C_OUTPUT_BRAM_106_DEPTH(C_OUTPUT_BRAM_106_DEPTH),
        .C_OUTPUT_BRAM_107_DEPTH(C_OUTPUT_BRAM_107_DEPTH),
        .C_OUTPUT_BRAM_108_DEPTH(C_OUTPUT_BRAM_108_DEPTH),
        .C_OUTPUT_BRAM_109_DEPTH(C_OUTPUT_BRAM_109_DEPTH),
        .C_OUTPUT_BRAM_110_DEPTH(C_OUTPUT_BRAM_110_DEPTH),
        .C_OUTPUT_BRAM_111_DEPTH(C_OUTPUT_BRAM_111_DEPTH),
        .C_OUTPUT_BRAM_112_DEPTH(C_OUTPUT_BRAM_112_DEPTH),
        .C_OUTPUT_BRAM_113_DEPTH(C_OUTPUT_BRAM_113_DEPTH),
        .C_OUTPUT_BRAM_114_DEPTH(C_OUTPUT_BRAM_114_DEPTH),
        .C_OUTPUT_BRAM_115_DEPTH(C_OUTPUT_BRAM_115_DEPTH),
        .C_OUTPUT_BRAM_116_DEPTH(C_OUTPUT_BRAM_116_DEPTH),
        .C_OUTPUT_BRAM_117_DEPTH(C_OUTPUT_BRAM_117_DEPTH),
        .C_OUTPUT_BRAM_118_DEPTH(C_OUTPUT_BRAM_118_DEPTH),
        .C_OUTPUT_BRAM_119_DEPTH(C_OUTPUT_BRAM_119_DEPTH),
        .C_OUTPUT_BRAM_120_DEPTH(C_OUTPUT_BRAM_120_DEPTH),
        .C_OUTPUT_BRAM_121_DEPTH(C_OUTPUT_BRAM_121_DEPTH),
        .C_OUTPUT_BRAM_122_DEPTH(C_OUTPUT_BRAM_122_DEPTH),
        .C_OUTPUT_BRAM_123_DEPTH(C_OUTPUT_BRAM_123_DEPTH),
        .C_OUTPUT_BRAM_124_DEPTH(C_OUTPUT_BRAM_124_DEPTH),
        .C_OUTPUT_BRAM_125_DEPTH(C_OUTPUT_BRAM_125_DEPTH),
        .C_OUTPUT_BRAM_126_DEPTH(C_OUTPUT_BRAM_126_DEPTH),
        .C_OUTPUT_BRAM_127_DEPTH(C_OUTPUT_BRAM_127_DEPTH),
        .C_OUTPUT_BRAM_0_DMWIDTH(C_OUTPUT_BRAM_0_DMWIDTH),
        .C_OUTPUT_BRAM_1_DMWIDTH(C_OUTPUT_BRAM_1_DMWIDTH),
        .C_OUTPUT_BRAM_2_DMWIDTH(C_OUTPUT_BRAM_2_DMWIDTH),
        .C_OUTPUT_BRAM_3_DMWIDTH(C_OUTPUT_BRAM_3_DMWIDTH),
        .C_OUTPUT_BRAM_4_DMWIDTH(C_OUTPUT_BRAM_4_DMWIDTH),
        .C_OUTPUT_BRAM_5_DMWIDTH(C_OUTPUT_BRAM_5_DMWIDTH),
        .C_OUTPUT_BRAM_6_DMWIDTH(C_OUTPUT_BRAM_6_DMWIDTH),
        .C_OUTPUT_BRAM_7_DMWIDTH(C_OUTPUT_BRAM_7_DMWIDTH),
        .C_OUTPUT_BRAM_8_DMWIDTH(C_OUTPUT_BRAM_8_DMWIDTH),
        .C_OUTPUT_BRAM_9_DMWIDTH(C_OUTPUT_BRAM_9_DMWIDTH),
        .C_OUTPUT_BRAM_10_DMWIDTH(C_OUTPUT_BRAM_10_DMWIDTH),
        .C_OUTPUT_BRAM_11_DMWIDTH(C_OUTPUT_BRAM_11_DMWIDTH),
        .C_OUTPUT_BRAM_12_DMWIDTH(C_OUTPUT_BRAM_12_DMWIDTH),
        .C_OUTPUT_BRAM_13_DMWIDTH(C_OUTPUT_BRAM_13_DMWIDTH),
        .C_OUTPUT_BRAM_14_DMWIDTH(C_OUTPUT_BRAM_14_DMWIDTH),
        .C_OUTPUT_BRAM_15_DMWIDTH(C_OUTPUT_BRAM_15_DMWIDTH),
        .C_OUTPUT_BRAM_16_DMWIDTH(C_OUTPUT_BRAM_16_DMWIDTH),
        .C_OUTPUT_BRAM_17_DMWIDTH(C_OUTPUT_BRAM_17_DMWIDTH),
        .C_OUTPUT_BRAM_18_DMWIDTH(C_OUTPUT_BRAM_18_DMWIDTH),
        .C_OUTPUT_BRAM_19_DMWIDTH(C_OUTPUT_BRAM_19_DMWIDTH),
        .C_OUTPUT_BRAM_20_DMWIDTH(C_OUTPUT_BRAM_20_DMWIDTH),
        .C_OUTPUT_BRAM_21_DMWIDTH(C_OUTPUT_BRAM_21_DMWIDTH),
        .C_OUTPUT_BRAM_22_DMWIDTH(C_OUTPUT_BRAM_22_DMWIDTH),
        .C_OUTPUT_BRAM_23_DMWIDTH(C_OUTPUT_BRAM_23_DMWIDTH),
        .C_OUTPUT_BRAM_24_DMWIDTH(C_OUTPUT_BRAM_24_DMWIDTH),
        .C_OUTPUT_BRAM_25_DMWIDTH(C_OUTPUT_BRAM_25_DMWIDTH),
        .C_OUTPUT_BRAM_26_DMWIDTH(C_OUTPUT_BRAM_26_DMWIDTH),
        .C_OUTPUT_BRAM_27_DMWIDTH(C_OUTPUT_BRAM_27_DMWIDTH),
        .C_OUTPUT_BRAM_28_DMWIDTH(C_OUTPUT_BRAM_28_DMWIDTH),
        .C_OUTPUT_BRAM_29_DMWIDTH(C_OUTPUT_BRAM_29_DMWIDTH),
        .C_OUTPUT_BRAM_30_DMWIDTH(C_OUTPUT_BRAM_30_DMWIDTH),
        .C_OUTPUT_BRAM_31_DMWIDTH(C_OUTPUT_BRAM_31_DMWIDTH),
        .C_OUTPUT_BRAM_32_DMWIDTH(C_OUTPUT_BRAM_32_DMWIDTH),
        .C_OUTPUT_BRAM_33_DMWIDTH(C_OUTPUT_BRAM_33_DMWIDTH),
        .C_OUTPUT_BRAM_34_DMWIDTH(C_OUTPUT_BRAM_34_DMWIDTH),
        .C_OUTPUT_BRAM_35_DMWIDTH(C_OUTPUT_BRAM_35_DMWIDTH),
        .C_OUTPUT_BRAM_36_DMWIDTH(C_OUTPUT_BRAM_36_DMWIDTH),
        .C_OUTPUT_BRAM_37_DMWIDTH(C_OUTPUT_BRAM_37_DMWIDTH),
        .C_OUTPUT_BRAM_38_DMWIDTH(C_OUTPUT_BRAM_38_DMWIDTH),
        .C_OUTPUT_BRAM_39_DMWIDTH(C_OUTPUT_BRAM_39_DMWIDTH),
        .C_OUTPUT_BRAM_40_DMWIDTH(C_OUTPUT_BRAM_40_DMWIDTH),
        .C_OUTPUT_BRAM_41_DMWIDTH(C_OUTPUT_BRAM_41_DMWIDTH),
        .C_OUTPUT_BRAM_42_DMWIDTH(C_OUTPUT_BRAM_42_DMWIDTH),
        .C_OUTPUT_BRAM_43_DMWIDTH(C_OUTPUT_BRAM_43_DMWIDTH),
        .C_OUTPUT_BRAM_44_DMWIDTH(C_OUTPUT_BRAM_44_DMWIDTH),
        .C_OUTPUT_BRAM_45_DMWIDTH(C_OUTPUT_BRAM_45_DMWIDTH),
        .C_OUTPUT_BRAM_46_DMWIDTH(C_OUTPUT_BRAM_46_DMWIDTH),
        .C_OUTPUT_BRAM_47_DMWIDTH(C_OUTPUT_BRAM_47_DMWIDTH),
        .C_OUTPUT_BRAM_48_DMWIDTH(C_OUTPUT_BRAM_48_DMWIDTH),
        .C_OUTPUT_BRAM_49_DMWIDTH(C_OUTPUT_BRAM_49_DMWIDTH),
        .C_OUTPUT_BRAM_50_DMWIDTH(C_OUTPUT_BRAM_50_DMWIDTH),
        .C_OUTPUT_BRAM_51_DMWIDTH(C_OUTPUT_BRAM_51_DMWIDTH),
        .C_OUTPUT_BRAM_52_DMWIDTH(C_OUTPUT_BRAM_52_DMWIDTH),
        .C_OUTPUT_BRAM_53_DMWIDTH(C_OUTPUT_BRAM_53_DMWIDTH),
        .C_OUTPUT_BRAM_54_DMWIDTH(C_OUTPUT_BRAM_54_DMWIDTH),
        .C_OUTPUT_BRAM_55_DMWIDTH(C_OUTPUT_BRAM_55_DMWIDTH),
        .C_OUTPUT_BRAM_56_DMWIDTH(C_OUTPUT_BRAM_56_DMWIDTH),
        .C_OUTPUT_BRAM_57_DMWIDTH(C_OUTPUT_BRAM_57_DMWIDTH),
        .C_OUTPUT_BRAM_58_DMWIDTH(C_OUTPUT_BRAM_58_DMWIDTH),
        .C_OUTPUT_BRAM_59_DMWIDTH(C_OUTPUT_BRAM_59_DMWIDTH),
        .C_OUTPUT_BRAM_60_DMWIDTH(C_OUTPUT_BRAM_60_DMWIDTH),
        .C_OUTPUT_BRAM_61_DMWIDTH(C_OUTPUT_BRAM_61_DMWIDTH),
        .C_OUTPUT_BRAM_62_DMWIDTH(C_OUTPUT_BRAM_62_DMWIDTH),
        .C_OUTPUT_BRAM_63_DMWIDTH(C_OUTPUT_BRAM_63_DMWIDTH),
        .C_OUTPUT_BRAM_64_DMWIDTH(C_OUTPUT_BRAM_64_DMWIDTH),
        .C_OUTPUT_BRAM_65_DMWIDTH(C_OUTPUT_BRAM_65_DMWIDTH),
        .C_OUTPUT_BRAM_66_DMWIDTH(C_OUTPUT_BRAM_66_DMWIDTH),
        .C_OUTPUT_BRAM_67_DMWIDTH(C_OUTPUT_BRAM_67_DMWIDTH),
        .C_OUTPUT_BRAM_68_DMWIDTH(C_OUTPUT_BRAM_68_DMWIDTH),
        .C_OUTPUT_BRAM_69_DMWIDTH(C_OUTPUT_BRAM_69_DMWIDTH),
        .C_OUTPUT_BRAM_70_DMWIDTH(C_OUTPUT_BRAM_70_DMWIDTH),
        .C_OUTPUT_BRAM_71_DMWIDTH(C_OUTPUT_BRAM_71_DMWIDTH),
        .C_OUTPUT_BRAM_72_DMWIDTH(C_OUTPUT_BRAM_72_DMWIDTH),
        .C_OUTPUT_BRAM_73_DMWIDTH(C_OUTPUT_BRAM_73_DMWIDTH),
        .C_OUTPUT_BRAM_74_DMWIDTH(C_OUTPUT_BRAM_74_DMWIDTH),
        .C_OUTPUT_BRAM_75_DMWIDTH(C_OUTPUT_BRAM_75_DMWIDTH),
        .C_OUTPUT_BRAM_76_DMWIDTH(C_OUTPUT_BRAM_76_DMWIDTH),
        .C_OUTPUT_BRAM_77_DMWIDTH(C_OUTPUT_BRAM_77_DMWIDTH),
        .C_OUTPUT_BRAM_78_DMWIDTH(C_OUTPUT_BRAM_78_DMWIDTH),
        .C_OUTPUT_BRAM_79_DMWIDTH(C_OUTPUT_BRAM_79_DMWIDTH),
        .C_OUTPUT_BRAM_80_DMWIDTH(C_OUTPUT_BRAM_80_DMWIDTH),
        .C_OUTPUT_BRAM_81_DMWIDTH(C_OUTPUT_BRAM_81_DMWIDTH),
        .C_OUTPUT_BRAM_82_DMWIDTH(C_OUTPUT_BRAM_82_DMWIDTH),
        .C_OUTPUT_BRAM_83_DMWIDTH(C_OUTPUT_BRAM_83_DMWIDTH),
        .C_OUTPUT_BRAM_84_DMWIDTH(C_OUTPUT_BRAM_84_DMWIDTH),
        .C_OUTPUT_BRAM_85_DMWIDTH(C_OUTPUT_BRAM_85_DMWIDTH),
        .C_OUTPUT_BRAM_86_DMWIDTH(C_OUTPUT_BRAM_86_DMWIDTH),
        .C_OUTPUT_BRAM_87_DMWIDTH(C_OUTPUT_BRAM_87_DMWIDTH),
        .C_OUTPUT_BRAM_88_DMWIDTH(C_OUTPUT_BRAM_88_DMWIDTH),
        .C_OUTPUT_BRAM_89_DMWIDTH(C_OUTPUT_BRAM_89_DMWIDTH),
        .C_OUTPUT_BRAM_90_DMWIDTH(C_OUTPUT_BRAM_90_DMWIDTH),
        .C_OUTPUT_BRAM_91_DMWIDTH(C_OUTPUT_BRAM_91_DMWIDTH),
        .C_OUTPUT_BRAM_92_DMWIDTH(C_OUTPUT_BRAM_92_DMWIDTH),
        .C_OUTPUT_BRAM_93_DMWIDTH(C_OUTPUT_BRAM_93_DMWIDTH),
        .C_OUTPUT_BRAM_94_DMWIDTH(C_OUTPUT_BRAM_94_DMWIDTH),
        .C_OUTPUT_BRAM_95_DMWIDTH(C_OUTPUT_BRAM_95_DMWIDTH),
        .C_OUTPUT_BRAM_96_DMWIDTH(C_OUTPUT_BRAM_96_DMWIDTH),
        .C_OUTPUT_BRAM_97_DMWIDTH(C_OUTPUT_BRAM_97_DMWIDTH),
        .C_OUTPUT_BRAM_98_DMWIDTH(C_OUTPUT_BRAM_98_DMWIDTH),
        .C_OUTPUT_BRAM_99_DMWIDTH(C_OUTPUT_BRAM_99_DMWIDTH),
        .C_OUTPUT_BRAM_100_DMWIDTH(C_OUTPUT_BRAM_100_DMWIDTH),
        .C_OUTPUT_BRAM_101_DMWIDTH(C_OUTPUT_BRAM_101_DMWIDTH),
        .C_OUTPUT_BRAM_102_DMWIDTH(C_OUTPUT_BRAM_102_DMWIDTH),
        .C_OUTPUT_BRAM_103_DMWIDTH(C_OUTPUT_BRAM_103_DMWIDTH),
        .C_OUTPUT_BRAM_104_DMWIDTH(C_OUTPUT_BRAM_104_DMWIDTH),
        .C_OUTPUT_BRAM_105_DMWIDTH(C_OUTPUT_BRAM_105_DMWIDTH),
        .C_OUTPUT_BRAM_106_DMWIDTH(C_OUTPUT_BRAM_106_DMWIDTH),
        .C_OUTPUT_BRAM_107_DMWIDTH(C_OUTPUT_BRAM_107_DMWIDTH),
        .C_OUTPUT_BRAM_108_DMWIDTH(C_OUTPUT_BRAM_108_DMWIDTH),
        .C_OUTPUT_BRAM_109_DMWIDTH(C_OUTPUT_BRAM_109_DMWIDTH),
        .C_OUTPUT_BRAM_110_DMWIDTH(C_OUTPUT_BRAM_110_DMWIDTH),
        .C_OUTPUT_BRAM_111_DMWIDTH(C_OUTPUT_BRAM_111_DMWIDTH),
        .C_OUTPUT_BRAM_112_DMWIDTH(C_OUTPUT_BRAM_112_DMWIDTH),
        .C_OUTPUT_BRAM_113_DMWIDTH(C_OUTPUT_BRAM_113_DMWIDTH),
        .C_OUTPUT_BRAM_114_DMWIDTH(C_OUTPUT_BRAM_114_DMWIDTH),
        .C_OUTPUT_BRAM_115_DMWIDTH(C_OUTPUT_BRAM_115_DMWIDTH),
        .C_OUTPUT_BRAM_116_DMWIDTH(C_OUTPUT_BRAM_116_DMWIDTH),
        .C_OUTPUT_BRAM_117_DMWIDTH(C_OUTPUT_BRAM_117_DMWIDTH),
        .C_OUTPUT_BRAM_118_DMWIDTH(C_OUTPUT_BRAM_118_DMWIDTH),
        .C_OUTPUT_BRAM_119_DMWIDTH(C_OUTPUT_BRAM_119_DMWIDTH),
        .C_OUTPUT_BRAM_120_DMWIDTH(C_OUTPUT_BRAM_120_DMWIDTH),
        .C_OUTPUT_BRAM_121_DMWIDTH(C_OUTPUT_BRAM_121_DMWIDTH),
        .C_OUTPUT_BRAM_122_DMWIDTH(C_OUTPUT_BRAM_122_DMWIDTH),
        .C_OUTPUT_BRAM_123_DMWIDTH(C_OUTPUT_BRAM_123_DMWIDTH),
        .C_OUTPUT_BRAM_124_DMWIDTH(C_OUTPUT_BRAM_124_DMWIDTH),
        .C_OUTPUT_BRAM_125_DMWIDTH(C_OUTPUT_BRAM_125_DMWIDTH),
        .C_OUTPUT_BRAM_126_DMWIDTH(C_OUTPUT_BRAM_126_DMWIDTH),
        .C_OUTPUT_BRAM_127_DMWIDTH(C_OUTPUT_BRAM_127_DMWIDTH),
        .C_OUTPUT_BRAM_0_MB_DEPTH(C_OUTPUT_BRAM_0_MB_DEPTH),
        .C_OUTPUT_BRAM_1_MB_DEPTH(C_OUTPUT_BRAM_1_MB_DEPTH),
        .C_OUTPUT_BRAM_2_MB_DEPTH(C_OUTPUT_BRAM_2_MB_DEPTH),
        .C_OUTPUT_BRAM_3_MB_DEPTH(C_OUTPUT_BRAM_3_MB_DEPTH),
        .C_OUTPUT_BRAM_4_MB_DEPTH(C_OUTPUT_BRAM_4_MB_DEPTH),
        .C_OUTPUT_BRAM_5_MB_DEPTH(C_OUTPUT_BRAM_5_MB_DEPTH),
        .C_OUTPUT_BRAM_6_MB_DEPTH(C_OUTPUT_BRAM_6_MB_DEPTH),
        .C_OUTPUT_BRAM_7_MB_DEPTH(C_OUTPUT_BRAM_7_MB_DEPTH),
        .C_OUTPUT_BRAM_8_MB_DEPTH(C_OUTPUT_BRAM_8_MB_DEPTH),
        .C_OUTPUT_BRAM_9_MB_DEPTH(C_OUTPUT_BRAM_9_MB_DEPTH),
        .C_OUTPUT_BRAM_10_MB_DEPTH(C_OUTPUT_BRAM_10_MB_DEPTH),
        .C_OUTPUT_BRAM_11_MB_DEPTH(C_OUTPUT_BRAM_11_MB_DEPTH),
        .C_OUTPUT_BRAM_12_MB_DEPTH(C_OUTPUT_BRAM_12_MB_DEPTH),
        .C_OUTPUT_BRAM_13_MB_DEPTH(C_OUTPUT_BRAM_13_MB_DEPTH),
        .C_OUTPUT_BRAM_14_MB_DEPTH(C_OUTPUT_BRAM_14_MB_DEPTH),
        .C_OUTPUT_BRAM_15_MB_DEPTH(C_OUTPUT_BRAM_15_MB_DEPTH),
        .C_OUTPUT_BRAM_16_MB_DEPTH(C_OUTPUT_BRAM_16_MB_DEPTH),
        .C_OUTPUT_BRAM_17_MB_DEPTH(C_OUTPUT_BRAM_17_MB_DEPTH),
        .C_OUTPUT_BRAM_18_MB_DEPTH(C_OUTPUT_BRAM_18_MB_DEPTH),
        .C_OUTPUT_BRAM_19_MB_DEPTH(C_OUTPUT_BRAM_19_MB_DEPTH),
        .C_OUTPUT_BRAM_20_MB_DEPTH(C_OUTPUT_BRAM_20_MB_DEPTH),
        .C_OUTPUT_BRAM_21_MB_DEPTH(C_OUTPUT_BRAM_21_MB_DEPTH),
        .C_OUTPUT_BRAM_22_MB_DEPTH(C_OUTPUT_BRAM_22_MB_DEPTH),
        .C_OUTPUT_BRAM_23_MB_DEPTH(C_OUTPUT_BRAM_23_MB_DEPTH),
        .C_OUTPUT_BRAM_24_MB_DEPTH(C_OUTPUT_BRAM_24_MB_DEPTH),
        .C_OUTPUT_BRAM_25_MB_DEPTH(C_OUTPUT_BRAM_25_MB_DEPTH),
        .C_OUTPUT_BRAM_26_MB_DEPTH(C_OUTPUT_BRAM_26_MB_DEPTH),
        .C_OUTPUT_BRAM_27_MB_DEPTH(C_OUTPUT_BRAM_27_MB_DEPTH),
        .C_OUTPUT_BRAM_28_MB_DEPTH(C_OUTPUT_BRAM_28_MB_DEPTH),
        .C_OUTPUT_BRAM_29_MB_DEPTH(C_OUTPUT_BRAM_29_MB_DEPTH),
        .C_OUTPUT_BRAM_30_MB_DEPTH(C_OUTPUT_BRAM_30_MB_DEPTH),
        .C_OUTPUT_BRAM_31_MB_DEPTH(C_OUTPUT_BRAM_31_MB_DEPTH),
        .C_OUTPUT_BRAM_32_MB_DEPTH(C_OUTPUT_BRAM_32_MB_DEPTH),
        .C_OUTPUT_BRAM_33_MB_DEPTH(C_OUTPUT_BRAM_33_MB_DEPTH),
        .C_OUTPUT_BRAM_34_MB_DEPTH(C_OUTPUT_BRAM_34_MB_DEPTH),
        .C_OUTPUT_BRAM_35_MB_DEPTH(C_OUTPUT_BRAM_35_MB_DEPTH),
        .C_OUTPUT_BRAM_36_MB_DEPTH(C_OUTPUT_BRAM_36_MB_DEPTH),
        .C_OUTPUT_BRAM_37_MB_DEPTH(C_OUTPUT_BRAM_37_MB_DEPTH),
        .C_OUTPUT_BRAM_38_MB_DEPTH(C_OUTPUT_BRAM_38_MB_DEPTH),
        .C_OUTPUT_BRAM_39_MB_DEPTH(C_OUTPUT_BRAM_39_MB_DEPTH),
        .C_OUTPUT_BRAM_40_MB_DEPTH(C_OUTPUT_BRAM_40_MB_DEPTH),
        .C_OUTPUT_BRAM_41_MB_DEPTH(C_OUTPUT_BRAM_41_MB_DEPTH),
        .C_OUTPUT_BRAM_42_MB_DEPTH(C_OUTPUT_BRAM_42_MB_DEPTH),
        .C_OUTPUT_BRAM_43_MB_DEPTH(C_OUTPUT_BRAM_43_MB_DEPTH),
        .C_OUTPUT_BRAM_44_MB_DEPTH(C_OUTPUT_BRAM_44_MB_DEPTH),
        .C_OUTPUT_BRAM_45_MB_DEPTH(C_OUTPUT_BRAM_45_MB_DEPTH),
        .C_OUTPUT_BRAM_46_MB_DEPTH(C_OUTPUT_BRAM_46_MB_DEPTH),
        .C_OUTPUT_BRAM_47_MB_DEPTH(C_OUTPUT_BRAM_47_MB_DEPTH),
        .C_OUTPUT_BRAM_48_MB_DEPTH(C_OUTPUT_BRAM_48_MB_DEPTH),
        .C_OUTPUT_BRAM_49_MB_DEPTH(C_OUTPUT_BRAM_49_MB_DEPTH),
        .C_OUTPUT_BRAM_50_MB_DEPTH(C_OUTPUT_BRAM_50_MB_DEPTH),
        .C_OUTPUT_BRAM_51_MB_DEPTH(C_OUTPUT_BRAM_51_MB_DEPTH),
        .C_OUTPUT_BRAM_52_MB_DEPTH(C_OUTPUT_BRAM_52_MB_DEPTH),
        .C_OUTPUT_BRAM_53_MB_DEPTH(C_OUTPUT_BRAM_53_MB_DEPTH),
        .C_OUTPUT_BRAM_54_MB_DEPTH(C_OUTPUT_BRAM_54_MB_DEPTH),
        .C_OUTPUT_BRAM_55_MB_DEPTH(C_OUTPUT_BRAM_55_MB_DEPTH),
        .C_OUTPUT_BRAM_56_MB_DEPTH(C_OUTPUT_BRAM_56_MB_DEPTH),
        .C_OUTPUT_BRAM_57_MB_DEPTH(C_OUTPUT_BRAM_57_MB_DEPTH),
        .C_OUTPUT_BRAM_58_MB_DEPTH(C_OUTPUT_BRAM_58_MB_DEPTH),
        .C_OUTPUT_BRAM_59_MB_DEPTH(C_OUTPUT_BRAM_59_MB_DEPTH),
        .C_OUTPUT_BRAM_60_MB_DEPTH(C_OUTPUT_BRAM_60_MB_DEPTH),
        .C_OUTPUT_BRAM_61_MB_DEPTH(C_OUTPUT_BRAM_61_MB_DEPTH),
        .C_OUTPUT_BRAM_62_MB_DEPTH(C_OUTPUT_BRAM_62_MB_DEPTH),
        .C_OUTPUT_BRAM_63_MB_DEPTH(C_OUTPUT_BRAM_63_MB_DEPTH),
        .C_OUTPUT_BRAM_64_MB_DEPTH(C_OUTPUT_BRAM_64_MB_DEPTH),
        .C_OUTPUT_BRAM_65_MB_DEPTH(C_OUTPUT_BRAM_65_MB_DEPTH),
        .C_OUTPUT_BRAM_66_MB_DEPTH(C_OUTPUT_BRAM_66_MB_DEPTH),
        .C_OUTPUT_BRAM_67_MB_DEPTH(C_OUTPUT_BRAM_67_MB_DEPTH),
        .C_OUTPUT_BRAM_68_MB_DEPTH(C_OUTPUT_BRAM_68_MB_DEPTH),
        .C_OUTPUT_BRAM_69_MB_DEPTH(C_OUTPUT_BRAM_69_MB_DEPTH),
        .C_OUTPUT_BRAM_70_MB_DEPTH(C_OUTPUT_BRAM_70_MB_DEPTH),
        .C_OUTPUT_BRAM_71_MB_DEPTH(C_OUTPUT_BRAM_71_MB_DEPTH),
        .C_OUTPUT_BRAM_72_MB_DEPTH(C_OUTPUT_BRAM_72_MB_DEPTH),
        .C_OUTPUT_BRAM_73_MB_DEPTH(C_OUTPUT_BRAM_73_MB_DEPTH),
        .C_OUTPUT_BRAM_74_MB_DEPTH(C_OUTPUT_BRAM_74_MB_DEPTH),
        .C_OUTPUT_BRAM_75_MB_DEPTH(C_OUTPUT_BRAM_75_MB_DEPTH),
        .C_OUTPUT_BRAM_76_MB_DEPTH(C_OUTPUT_BRAM_76_MB_DEPTH),
        .C_OUTPUT_BRAM_77_MB_DEPTH(C_OUTPUT_BRAM_77_MB_DEPTH),
        .C_OUTPUT_BRAM_78_MB_DEPTH(C_OUTPUT_BRAM_78_MB_DEPTH),
        .C_OUTPUT_BRAM_79_MB_DEPTH(C_OUTPUT_BRAM_79_MB_DEPTH),
        .C_OUTPUT_BRAM_80_MB_DEPTH(C_OUTPUT_BRAM_80_MB_DEPTH),
        .C_OUTPUT_BRAM_81_MB_DEPTH(C_OUTPUT_BRAM_81_MB_DEPTH),
        .C_OUTPUT_BRAM_82_MB_DEPTH(C_OUTPUT_BRAM_82_MB_DEPTH),
        .C_OUTPUT_BRAM_83_MB_DEPTH(C_OUTPUT_BRAM_83_MB_DEPTH),
        .C_OUTPUT_BRAM_84_MB_DEPTH(C_OUTPUT_BRAM_84_MB_DEPTH),
        .C_OUTPUT_BRAM_85_MB_DEPTH(C_OUTPUT_BRAM_85_MB_DEPTH),
        .C_OUTPUT_BRAM_86_MB_DEPTH(C_OUTPUT_BRAM_86_MB_DEPTH),
        .C_OUTPUT_BRAM_87_MB_DEPTH(C_OUTPUT_BRAM_87_MB_DEPTH),
        .C_OUTPUT_BRAM_88_MB_DEPTH(C_OUTPUT_BRAM_88_MB_DEPTH),
        .C_OUTPUT_BRAM_89_MB_DEPTH(C_OUTPUT_BRAM_89_MB_DEPTH),
        .C_OUTPUT_BRAM_90_MB_DEPTH(C_OUTPUT_BRAM_90_MB_DEPTH),
        .C_OUTPUT_BRAM_91_MB_DEPTH(C_OUTPUT_BRAM_91_MB_DEPTH),
        .C_OUTPUT_BRAM_92_MB_DEPTH(C_OUTPUT_BRAM_92_MB_DEPTH),
        .C_OUTPUT_BRAM_93_MB_DEPTH(C_OUTPUT_BRAM_93_MB_DEPTH),
        .C_OUTPUT_BRAM_94_MB_DEPTH(C_OUTPUT_BRAM_94_MB_DEPTH),
        .C_OUTPUT_BRAM_95_MB_DEPTH(C_OUTPUT_BRAM_95_MB_DEPTH),
        .C_OUTPUT_BRAM_96_MB_DEPTH(C_OUTPUT_BRAM_96_MB_DEPTH),
        .C_OUTPUT_BRAM_97_MB_DEPTH(C_OUTPUT_BRAM_97_MB_DEPTH),
        .C_OUTPUT_BRAM_98_MB_DEPTH(C_OUTPUT_BRAM_98_MB_DEPTH),
        .C_OUTPUT_BRAM_99_MB_DEPTH(C_OUTPUT_BRAM_99_MB_DEPTH),
        .C_OUTPUT_BRAM_100_MB_DEPTH(C_OUTPUT_BRAM_100_MB_DEPTH),
        .C_OUTPUT_BRAM_101_MB_DEPTH(C_OUTPUT_BRAM_101_MB_DEPTH),
        .C_OUTPUT_BRAM_102_MB_DEPTH(C_OUTPUT_BRAM_102_MB_DEPTH),
        .C_OUTPUT_BRAM_103_MB_DEPTH(C_OUTPUT_BRAM_103_MB_DEPTH),
        .C_OUTPUT_BRAM_104_MB_DEPTH(C_OUTPUT_BRAM_104_MB_DEPTH),
        .C_OUTPUT_BRAM_105_MB_DEPTH(C_OUTPUT_BRAM_105_MB_DEPTH),
        .C_OUTPUT_BRAM_106_MB_DEPTH(C_OUTPUT_BRAM_106_MB_DEPTH),
        .C_OUTPUT_BRAM_107_MB_DEPTH(C_OUTPUT_BRAM_107_MB_DEPTH),
        .C_OUTPUT_BRAM_108_MB_DEPTH(C_OUTPUT_BRAM_108_MB_DEPTH),
        .C_OUTPUT_BRAM_109_MB_DEPTH(C_OUTPUT_BRAM_109_MB_DEPTH),
        .C_OUTPUT_BRAM_110_MB_DEPTH(C_OUTPUT_BRAM_110_MB_DEPTH),
        .C_OUTPUT_BRAM_111_MB_DEPTH(C_OUTPUT_BRAM_111_MB_DEPTH),
        .C_OUTPUT_BRAM_112_MB_DEPTH(C_OUTPUT_BRAM_112_MB_DEPTH),
        .C_OUTPUT_BRAM_113_MB_DEPTH(C_OUTPUT_BRAM_113_MB_DEPTH),
        .C_OUTPUT_BRAM_114_MB_DEPTH(C_OUTPUT_BRAM_114_MB_DEPTH),
        .C_OUTPUT_BRAM_115_MB_DEPTH(C_OUTPUT_BRAM_115_MB_DEPTH),
        .C_OUTPUT_BRAM_116_MB_DEPTH(C_OUTPUT_BRAM_116_MB_DEPTH),
        .C_OUTPUT_BRAM_117_MB_DEPTH(C_OUTPUT_BRAM_117_MB_DEPTH),
        .C_OUTPUT_BRAM_118_MB_DEPTH(C_OUTPUT_BRAM_118_MB_DEPTH),
        .C_OUTPUT_BRAM_119_MB_DEPTH(C_OUTPUT_BRAM_119_MB_DEPTH),
        .C_OUTPUT_BRAM_120_MB_DEPTH(C_OUTPUT_BRAM_120_MB_DEPTH),
        .C_OUTPUT_BRAM_121_MB_DEPTH(C_OUTPUT_BRAM_121_MB_DEPTH),
        .C_OUTPUT_BRAM_122_MB_DEPTH(C_OUTPUT_BRAM_122_MB_DEPTH),
        .C_OUTPUT_BRAM_123_MB_DEPTH(C_OUTPUT_BRAM_123_MB_DEPTH),
        .C_OUTPUT_BRAM_124_MB_DEPTH(C_OUTPUT_BRAM_124_MB_DEPTH),
        .C_OUTPUT_BRAM_125_MB_DEPTH(C_OUTPUT_BRAM_125_MB_DEPTH),
        .C_OUTPUT_BRAM_126_MB_DEPTH(C_OUTPUT_BRAM_126_MB_DEPTH),
        .C_OUTPUT_BRAM_127_MB_DEPTH(C_OUTPUT_BRAM_127_MB_DEPTH),
        .C_OUTPUT_BRAM_0_ADDR_WIDTH(C_OUTPUT_BRAM_0_ADDR_WIDTH),
        .C_OUTPUT_BRAM_1_ADDR_WIDTH(C_OUTPUT_BRAM_1_ADDR_WIDTH),
        .C_OUTPUT_BRAM_2_ADDR_WIDTH(C_OUTPUT_BRAM_2_ADDR_WIDTH),
        .C_OUTPUT_BRAM_3_ADDR_WIDTH(C_OUTPUT_BRAM_3_ADDR_WIDTH),
        .C_OUTPUT_BRAM_4_ADDR_WIDTH(C_OUTPUT_BRAM_4_ADDR_WIDTH),
        .C_OUTPUT_BRAM_5_ADDR_WIDTH(C_OUTPUT_BRAM_5_ADDR_WIDTH),
        .C_OUTPUT_BRAM_6_ADDR_WIDTH(C_OUTPUT_BRAM_6_ADDR_WIDTH),
        .C_OUTPUT_BRAM_7_ADDR_WIDTH(C_OUTPUT_BRAM_7_ADDR_WIDTH),
        .C_OUTPUT_BRAM_8_ADDR_WIDTH(C_OUTPUT_BRAM_8_ADDR_WIDTH),
        .C_OUTPUT_BRAM_9_ADDR_WIDTH(C_OUTPUT_BRAM_9_ADDR_WIDTH),
        .C_OUTPUT_BRAM_10_ADDR_WIDTH(C_OUTPUT_BRAM_10_ADDR_WIDTH),
        .C_OUTPUT_BRAM_11_ADDR_WIDTH(C_OUTPUT_BRAM_11_ADDR_WIDTH),
        .C_OUTPUT_BRAM_12_ADDR_WIDTH(C_OUTPUT_BRAM_12_ADDR_WIDTH),
        .C_OUTPUT_BRAM_13_ADDR_WIDTH(C_OUTPUT_BRAM_13_ADDR_WIDTH),
        .C_OUTPUT_BRAM_14_ADDR_WIDTH(C_OUTPUT_BRAM_14_ADDR_WIDTH),
        .C_OUTPUT_BRAM_15_ADDR_WIDTH(C_OUTPUT_BRAM_15_ADDR_WIDTH),
        .C_OUTPUT_BRAM_16_ADDR_WIDTH(C_OUTPUT_BRAM_16_ADDR_WIDTH),
        .C_OUTPUT_BRAM_17_ADDR_WIDTH(C_OUTPUT_BRAM_17_ADDR_WIDTH),
        .C_OUTPUT_BRAM_18_ADDR_WIDTH(C_OUTPUT_BRAM_18_ADDR_WIDTH),
        .C_OUTPUT_BRAM_19_ADDR_WIDTH(C_OUTPUT_BRAM_19_ADDR_WIDTH),
        .C_OUTPUT_BRAM_20_ADDR_WIDTH(C_OUTPUT_BRAM_20_ADDR_WIDTH),
        .C_OUTPUT_BRAM_21_ADDR_WIDTH(C_OUTPUT_BRAM_21_ADDR_WIDTH),
        .C_OUTPUT_BRAM_22_ADDR_WIDTH(C_OUTPUT_BRAM_22_ADDR_WIDTH),
        .C_OUTPUT_BRAM_23_ADDR_WIDTH(C_OUTPUT_BRAM_23_ADDR_WIDTH),
        .C_OUTPUT_BRAM_24_ADDR_WIDTH(C_OUTPUT_BRAM_24_ADDR_WIDTH),
        .C_OUTPUT_BRAM_25_ADDR_WIDTH(C_OUTPUT_BRAM_25_ADDR_WIDTH),
        .C_OUTPUT_BRAM_26_ADDR_WIDTH(C_OUTPUT_BRAM_26_ADDR_WIDTH),
        .C_OUTPUT_BRAM_27_ADDR_WIDTH(C_OUTPUT_BRAM_27_ADDR_WIDTH),
        .C_OUTPUT_BRAM_28_ADDR_WIDTH(C_OUTPUT_BRAM_28_ADDR_WIDTH),
        .C_OUTPUT_BRAM_29_ADDR_WIDTH(C_OUTPUT_BRAM_29_ADDR_WIDTH),
        .C_OUTPUT_BRAM_30_ADDR_WIDTH(C_OUTPUT_BRAM_30_ADDR_WIDTH),
        .C_OUTPUT_BRAM_31_ADDR_WIDTH(C_OUTPUT_BRAM_31_ADDR_WIDTH),
        .C_OUTPUT_BRAM_32_ADDR_WIDTH(C_OUTPUT_BRAM_32_ADDR_WIDTH),
        .C_OUTPUT_BRAM_33_ADDR_WIDTH(C_OUTPUT_BRAM_33_ADDR_WIDTH),
        .C_OUTPUT_BRAM_34_ADDR_WIDTH(C_OUTPUT_BRAM_34_ADDR_WIDTH),
        .C_OUTPUT_BRAM_35_ADDR_WIDTH(C_OUTPUT_BRAM_35_ADDR_WIDTH),
        .C_OUTPUT_BRAM_36_ADDR_WIDTH(C_OUTPUT_BRAM_36_ADDR_WIDTH),
        .C_OUTPUT_BRAM_37_ADDR_WIDTH(C_OUTPUT_BRAM_37_ADDR_WIDTH),
        .C_OUTPUT_BRAM_38_ADDR_WIDTH(C_OUTPUT_BRAM_38_ADDR_WIDTH),
        .C_OUTPUT_BRAM_39_ADDR_WIDTH(C_OUTPUT_BRAM_39_ADDR_WIDTH),
        .C_OUTPUT_BRAM_40_ADDR_WIDTH(C_OUTPUT_BRAM_40_ADDR_WIDTH),
        .C_OUTPUT_BRAM_41_ADDR_WIDTH(C_OUTPUT_BRAM_41_ADDR_WIDTH),
        .C_OUTPUT_BRAM_42_ADDR_WIDTH(C_OUTPUT_BRAM_42_ADDR_WIDTH),
        .C_OUTPUT_BRAM_43_ADDR_WIDTH(C_OUTPUT_BRAM_43_ADDR_WIDTH),
        .C_OUTPUT_BRAM_44_ADDR_WIDTH(C_OUTPUT_BRAM_44_ADDR_WIDTH),
        .C_OUTPUT_BRAM_45_ADDR_WIDTH(C_OUTPUT_BRAM_45_ADDR_WIDTH),
        .C_OUTPUT_BRAM_46_ADDR_WIDTH(C_OUTPUT_BRAM_46_ADDR_WIDTH),
        .C_OUTPUT_BRAM_47_ADDR_WIDTH(C_OUTPUT_BRAM_47_ADDR_WIDTH),
        .C_OUTPUT_BRAM_48_ADDR_WIDTH(C_OUTPUT_BRAM_48_ADDR_WIDTH),
        .C_OUTPUT_BRAM_49_ADDR_WIDTH(C_OUTPUT_BRAM_49_ADDR_WIDTH),
        .C_OUTPUT_BRAM_50_ADDR_WIDTH(C_OUTPUT_BRAM_50_ADDR_WIDTH),
        .C_OUTPUT_BRAM_51_ADDR_WIDTH(C_OUTPUT_BRAM_51_ADDR_WIDTH),
        .C_OUTPUT_BRAM_52_ADDR_WIDTH(C_OUTPUT_BRAM_52_ADDR_WIDTH),
        .C_OUTPUT_BRAM_53_ADDR_WIDTH(C_OUTPUT_BRAM_53_ADDR_WIDTH),
        .C_OUTPUT_BRAM_54_ADDR_WIDTH(C_OUTPUT_BRAM_54_ADDR_WIDTH),
        .C_OUTPUT_BRAM_55_ADDR_WIDTH(C_OUTPUT_BRAM_55_ADDR_WIDTH),
        .C_OUTPUT_BRAM_56_ADDR_WIDTH(C_OUTPUT_BRAM_56_ADDR_WIDTH),
        .C_OUTPUT_BRAM_57_ADDR_WIDTH(C_OUTPUT_BRAM_57_ADDR_WIDTH),
        .C_OUTPUT_BRAM_58_ADDR_WIDTH(C_OUTPUT_BRAM_58_ADDR_WIDTH),
        .C_OUTPUT_BRAM_59_ADDR_WIDTH(C_OUTPUT_BRAM_59_ADDR_WIDTH),
        .C_OUTPUT_BRAM_60_ADDR_WIDTH(C_OUTPUT_BRAM_60_ADDR_WIDTH),
        .C_OUTPUT_BRAM_61_ADDR_WIDTH(C_OUTPUT_BRAM_61_ADDR_WIDTH),
        .C_OUTPUT_BRAM_62_ADDR_WIDTH(C_OUTPUT_BRAM_62_ADDR_WIDTH),
        .C_OUTPUT_BRAM_63_ADDR_WIDTH(C_OUTPUT_BRAM_63_ADDR_WIDTH),
        .C_OUTPUT_BRAM_64_ADDR_WIDTH(C_OUTPUT_BRAM_64_ADDR_WIDTH),
        .C_OUTPUT_BRAM_65_ADDR_WIDTH(C_OUTPUT_BRAM_65_ADDR_WIDTH),
        .C_OUTPUT_BRAM_66_ADDR_WIDTH(C_OUTPUT_BRAM_66_ADDR_WIDTH),
        .C_OUTPUT_BRAM_67_ADDR_WIDTH(C_OUTPUT_BRAM_67_ADDR_WIDTH),
        .C_OUTPUT_BRAM_68_ADDR_WIDTH(C_OUTPUT_BRAM_68_ADDR_WIDTH),
        .C_OUTPUT_BRAM_69_ADDR_WIDTH(C_OUTPUT_BRAM_69_ADDR_WIDTH),
        .C_OUTPUT_BRAM_70_ADDR_WIDTH(C_OUTPUT_BRAM_70_ADDR_WIDTH),
        .C_OUTPUT_BRAM_71_ADDR_WIDTH(C_OUTPUT_BRAM_71_ADDR_WIDTH),
        .C_OUTPUT_BRAM_72_ADDR_WIDTH(C_OUTPUT_BRAM_72_ADDR_WIDTH),
        .C_OUTPUT_BRAM_73_ADDR_WIDTH(C_OUTPUT_BRAM_73_ADDR_WIDTH),
        .C_OUTPUT_BRAM_74_ADDR_WIDTH(C_OUTPUT_BRAM_74_ADDR_WIDTH),
        .C_OUTPUT_BRAM_75_ADDR_WIDTH(C_OUTPUT_BRAM_75_ADDR_WIDTH),
        .C_OUTPUT_BRAM_76_ADDR_WIDTH(C_OUTPUT_BRAM_76_ADDR_WIDTH),
        .C_OUTPUT_BRAM_77_ADDR_WIDTH(C_OUTPUT_BRAM_77_ADDR_WIDTH),
        .C_OUTPUT_BRAM_78_ADDR_WIDTH(C_OUTPUT_BRAM_78_ADDR_WIDTH),
        .C_OUTPUT_BRAM_79_ADDR_WIDTH(C_OUTPUT_BRAM_79_ADDR_WIDTH),
        .C_OUTPUT_BRAM_80_ADDR_WIDTH(C_OUTPUT_BRAM_80_ADDR_WIDTH),
        .C_OUTPUT_BRAM_81_ADDR_WIDTH(C_OUTPUT_BRAM_81_ADDR_WIDTH),
        .C_OUTPUT_BRAM_82_ADDR_WIDTH(C_OUTPUT_BRAM_82_ADDR_WIDTH),
        .C_OUTPUT_BRAM_83_ADDR_WIDTH(C_OUTPUT_BRAM_83_ADDR_WIDTH),
        .C_OUTPUT_BRAM_84_ADDR_WIDTH(C_OUTPUT_BRAM_84_ADDR_WIDTH),
        .C_OUTPUT_BRAM_85_ADDR_WIDTH(C_OUTPUT_BRAM_85_ADDR_WIDTH),
        .C_OUTPUT_BRAM_86_ADDR_WIDTH(C_OUTPUT_BRAM_86_ADDR_WIDTH),
        .C_OUTPUT_BRAM_87_ADDR_WIDTH(C_OUTPUT_BRAM_87_ADDR_WIDTH),
        .C_OUTPUT_BRAM_88_ADDR_WIDTH(C_OUTPUT_BRAM_88_ADDR_WIDTH),
        .C_OUTPUT_BRAM_89_ADDR_WIDTH(C_OUTPUT_BRAM_89_ADDR_WIDTH),
        .C_OUTPUT_BRAM_90_ADDR_WIDTH(C_OUTPUT_BRAM_90_ADDR_WIDTH),
        .C_OUTPUT_BRAM_91_ADDR_WIDTH(C_OUTPUT_BRAM_91_ADDR_WIDTH),
        .C_OUTPUT_BRAM_92_ADDR_WIDTH(C_OUTPUT_BRAM_92_ADDR_WIDTH),
        .C_OUTPUT_BRAM_93_ADDR_WIDTH(C_OUTPUT_BRAM_93_ADDR_WIDTH),
        .C_OUTPUT_BRAM_94_ADDR_WIDTH(C_OUTPUT_BRAM_94_ADDR_WIDTH),
        .C_OUTPUT_BRAM_95_ADDR_WIDTH(C_OUTPUT_BRAM_95_ADDR_WIDTH),
        .C_OUTPUT_BRAM_96_ADDR_WIDTH(C_OUTPUT_BRAM_96_ADDR_WIDTH),
        .C_OUTPUT_BRAM_97_ADDR_WIDTH(C_OUTPUT_BRAM_97_ADDR_WIDTH),
        .C_OUTPUT_BRAM_98_ADDR_WIDTH(C_OUTPUT_BRAM_98_ADDR_WIDTH),
        .C_OUTPUT_BRAM_99_ADDR_WIDTH(C_OUTPUT_BRAM_99_ADDR_WIDTH),
        .C_OUTPUT_BRAM_100_ADDR_WIDTH(C_OUTPUT_BRAM_100_ADDR_WIDTH),
        .C_OUTPUT_BRAM_101_ADDR_WIDTH(C_OUTPUT_BRAM_101_ADDR_WIDTH),
        .C_OUTPUT_BRAM_102_ADDR_WIDTH(C_OUTPUT_BRAM_102_ADDR_WIDTH),
        .C_OUTPUT_BRAM_103_ADDR_WIDTH(C_OUTPUT_BRAM_103_ADDR_WIDTH),
        .C_OUTPUT_BRAM_104_ADDR_WIDTH(C_OUTPUT_BRAM_104_ADDR_WIDTH),
        .C_OUTPUT_BRAM_105_ADDR_WIDTH(C_OUTPUT_BRAM_105_ADDR_WIDTH),
        .C_OUTPUT_BRAM_106_ADDR_WIDTH(C_OUTPUT_BRAM_106_ADDR_WIDTH),
        .C_OUTPUT_BRAM_107_ADDR_WIDTH(C_OUTPUT_BRAM_107_ADDR_WIDTH),
        .C_OUTPUT_BRAM_108_ADDR_WIDTH(C_OUTPUT_BRAM_108_ADDR_WIDTH),
        .C_OUTPUT_BRAM_109_ADDR_WIDTH(C_OUTPUT_BRAM_109_ADDR_WIDTH),
        .C_OUTPUT_BRAM_110_ADDR_WIDTH(C_OUTPUT_BRAM_110_ADDR_WIDTH),
        .C_OUTPUT_BRAM_111_ADDR_WIDTH(C_OUTPUT_BRAM_111_ADDR_WIDTH),
        .C_OUTPUT_BRAM_112_ADDR_WIDTH(C_OUTPUT_BRAM_112_ADDR_WIDTH),
        .C_OUTPUT_BRAM_113_ADDR_WIDTH(C_OUTPUT_BRAM_113_ADDR_WIDTH),
        .C_OUTPUT_BRAM_114_ADDR_WIDTH(C_OUTPUT_BRAM_114_ADDR_WIDTH),
        .C_OUTPUT_BRAM_115_ADDR_WIDTH(C_OUTPUT_BRAM_115_ADDR_WIDTH),
        .C_OUTPUT_BRAM_116_ADDR_WIDTH(C_OUTPUT_BRAM_116_ADDR_WIDTH),
        .C_OUTPUT_BRAM_117_ADDR_WIDTH(C_OUTPUT_BRAM_117_ADDR_WIDTH),
        .C_OUTPUT_BRAM_118_ADDR_WIDTH(C_OUTPUT_BRAM_118_ADDR_WIDTH),
        .C_OUTPUT_BRAM_119_ADDR_WIDTH(C_OUTPUT_BRAM_119_ADDR_WIDTH),
        .C_OUTPUT_BRAM_120_ADDR_WIDTH(C_OUTPUT_BRAM_120_ADDR_WIDTH),
        .C_OUTPUT_BRAM_121_ADDR_WIDTH(C_OUTPUT_BRAM_121_ADDR_WIDTH),
        .C_OUTPUT_BRAM_122_ADDR_WIDTH(C_OUTPUT_BRAM_122_ADDR_WIDTH),
        .C_OUTPUT_BRAM_123_ADDR_WIDTH(C_OUTPUT_BRAM_123_ADDR_WIDTH),
        .C_OUTPUT_BRAM_124_ADDR_WIDTH(C_OUTPUT_BRAM_124_ADDR_WIDTH),
        .C_OUTPUT_BRAM_125_ADDR_WIDTH(C_OUTPUT_BRAM_125_ADDR_WIDTH),
        .C_OUTPUT_BRAM_126_ADDR_WIDTH(C_OUTPUT_BRAM_126_ADDR_WIDTH),
        .C_OUTPUT_BRAM_127_ADDR_WIDTH(C_OUTPUT_BRAM_127_ADDR_WIDTH)
    ) out_bram_args_i (
        .acc_clk(aclk),
        .dm_clk(s_axi_aclk),
        .aresetn(s_axi_aresetn),
        .acc_rstn(resetn),
        .outbram_allow(outbram_ctrl_allow),
        .acc_start(ap_start_single),
        .acc_done(ap_done),
        .outbram_ready(outbram_ctrl_ready),
        .outbram_canstart(outbram_ctrl_canstart),
        .outbram_depth(outbram_depth),
        .outbram_depth_write(outbram_depth_write),
        .m_axis_bram_0_tlast(m_axis_bram_0_tlast),
        .m_axis_bram_0_tvalid(m_axis_bram_0_tvalid),
        .m_axis_bram_0_tkeep(m_axis_bram_0_tkeep),
        .m_axis_bram_0_tstrb(m_axis_bram_0_tstrb),
        .m_axis_bram_0_tdata(m_axis_bram_0_tdata),
        .m_axis_bram_0_tready(m_axis_bram_0_tready),
        .ap_bram_0_addr0(ap_bram_oarg_0_addr0),
        .ap_bram_0_din0(ap_bram_oarg_0_din0),
        .ap_bram_0_dout0(ap_bram_oarg_0_dout0),
        .ap_bram_0_we0(ap_bram_oarg_0_we0),
        .ap_bram_0_en0(ap_bram_oarg_0_en0),
        .ap_bram_0_addr1(ap_bram_oarg_0_addr1),
        .ap_bram_0_din1(ap_bram_oarg_0_din1),
        .ap_bram_0_dout1(ap_bram_oarg_0_dout1),
        .ap_bram_0_we1(ap_bram_oarg_0_we1),
        .ap_bram_0_en1(ap_bram_oarg_0_en1),
        .m_axis_bram_1_tlast(m_axis_bram_1_tlast),
        .m_axis_bram_1_tvalid(m_axis_bram_1_tvalid),
        .m_axis_bram_1_tkeep(m_axis_bram_1_tkeep),
        .m_axis_bram_1_tstrb(m_axis_bram_1_tstrb),
        .m_axis_bram_1_tdata(m_axis_bram_1_tdata),
        .m_axis_bram_1_tready(m_axis_bram_1_tready),
        .ap_bram_1_addr0(ap_bram_oarg_1_addr0),
        .ap_bram_1_din0(ap_bram_oarg_1_din0),
        .ap_bram_1_dout0(ap_bram_oarg_1_dout0),
        .ap_bram_1_we0(ap_bram_oarg_1_we0),
        .ap_bram_1_en0(ap_bram_oarg_1_en0),
        .ap_bram_1_addr1(ap_bram_oarg_1_addr1),
        .ap_bram_1_din1(ap_bram_oarg_1_din1),
        .ap_bram_1_dout1(ap_bram_oarg_1_dout1),
        .ap_bram_1_we1(ap_bram_oarg_1_we1),
        .ap_bram_1_en1(ap_bram_oarg_1_en1),
        .m_axis_bram_2_tlast(m_axis_bram_2_tlast),
        .m_axis_bram_2_tvalid(m_axis_bram_2_tvalid),
        .m_axis_bram_2_tkeep(m_axis_bram_2_tkeep),
        .m_axis_bram_2_tstrb(m_axis_bram_2_tstrb),
        .m_axis_bram_2_tdata(m_axis_bram_2_tdata),
        .m_axis_bram_2_tready(m_axis_bram_2_tready),
        .ap_bram_2_addr0(ap_bram_oarg_2_addr0),
        .ap_bram_2_din0(ap_bram_oarg_2_din0),
        .ap_bram_2_dout0(ap_bram_oarg_2_dout0),
        .ap_bram_2_we0(ap_bram_oarg_2_we0),
        .ap_bram_2_en0(ap_bram_oarg_2_en0),
        .ap_bram_2_addr1(ap_bram_oarg_2_addr1),
        .ap_bram_2_din1(ap_bram_oarg_2_din1),
        .ap_bram_2_dout1(ap_bram_oarg_2_dout1),
        .ap_bram_2_we1(ap_bram_oarg_2_we1),
        .ap_bram_2_en1(ap_bram_oarg_2_en1),
        .m_axis_bram_3_tlast(m_axis_bram_3_tlast),
        .m_axis_bram_3_tvalid(m_axis_bram_3_tvalid),
        .m_axis_bram_3_tkeep(m_axis_bram_3_tkeep),
        .m_axis_bram_3_tstrb(m_axis_bram_3_tstrb),
        .m_axis_bram_3_tdata(m_axis_bram_3_tdata),
        .m_axis_bram_3_tready(m_axis_bram_3_tready),
        .ap_bram_3_addr0(ap_bram_oarg_3_addr0),
        .ap_bram_3_din0(ap_bram_oarg_3_din0),
        .ap_bram_3_dout0(ap_bram_oarg_3_dout0),
        .ap_bram_3_we0(ap_bram_oarg_3_we0),
        .ap_bram_3_en0(ap_bram_oarg_3_en0),
        .ap_bram_3_addr1(ap_bram_oarg_3_addr1),
        .ap_bram_3_din1(ap_bram_oarg_3_din1),
        .ap_bram_3_dout1(ap_bram_oarg_3_dout1),
        .ap_bram_3_we1(ap_bram_oarg_3_we1),
        .ap_bram_3_en1(ap_bram_oarg_3_en1),
        .m_axis_bram_4_tlast(m_axis_bram_4_tlast),
        .m_axis_bram_4_tvalid(m_axis_bram_4_tvalid),
        .m_axis_bram_4_tkeep(m_axis_bram_4_tkeep),
        .m_axis_bram_4_tstrb(m_axis_bram_4_tstrb),
        .m_axis_bram_4_tdata(m_axis_bram_4_tdata),
        .m_axis_bram_4_tready(m_axis_bram_4_tready),
        .ap_bram_4_addr0(ap_bram_oarg_4_addr0),
        .ap_bram_4_din0(ap_bram_oarg_4_din0),
        .ap_bram_4_dout0(ap_bram_oarg_4_dout0),
        .ap_bram_4_we0(ap_bram_oarg_4_we0),
        .ap_bram_4_en0(ap_bram_oarg_4_en0),
        .ap_bram_4_addr1(ap_bram_oarg_4_addr1),
        .ap_bram_4_din1(ap_bram_oarg_4_din1),
        .ap_bram_4_dout1(ap_bram_oarg_4_dout1),
        .ap_bram_4_we1(ap_bram_oarg_4_we1),
        .ap_bram_4_en1(ap_bram_oarg_4_en1),
        .m_axis_bram_5_tlast(m_axis_bram_5_tlast),
        .m_axis_bram_5_tvalid(m_axis_bram_5_tvalid),
        .m_axis_bram_5_tkeep(m_axis_bram_5_tkeep),
        .m_axis_bram_5_tstrb(m_axis_bram_5_tstrb),
        .m_axis_bram_5_tdata(m_axis_bram_5_tdata),
        .m_axis_bram_5_tready(m_axis_bram_5_tready),
        .ap_bram_5_addr0(ap_bram_oarg_5_addr0),
        .ap_bram_5_din0(ap_bram_oarg_5_din0),
        .ap_bram_5_dout0(ap_bram_oarg_5_dout0),
        .ap_bram_5_we0(ap_bram_oarg_5_we0),
        .ap_bram_5_en0(ap_bram_oarg_5_en0),
        .ap_bram_5_addr1(ap_bram_oarg_5_addr1),
        .ap_bram_5_din1(ap_bram_oarg_5_din1),
        .ap_bram_5_dout1(ap_bram_oarg_5_dout1),
        .ap_bram_5_we1(ap_bram_oarg_5_we1),
        .ap_bram_5_en1(ap_bram_oarg_5_en1),
        .m_axis_bram_6_tlast(m_axis_bram_6_tlast),
        .m_axis_bram_6_tvalid(m_axis_bram_6_tvalid),
        .m_axis_bram_6_tkeep(m_axis_bram_6_tkeep),
        .m_axis_bram_6_tstrb(m_axis_bram_6_tstrb),
        .m_axis_bram_6_tdata(m_axis_bram_6_tdata),
        .m_axis_bram_6_tready(m_axis_bram_6_tready),
        .ap_bram_6_addr0(ap_bram_oarg_6_addr0),
        .ap_bram_6_din0(ap_bram_oarg_6_din0),
        .ap_bram_6_dout0(ap_bram_oarg_6_dout0),
        .ap_bram_6_we0(ap_bram_oarg_6_we0),
        .ap_bram_6_en0(ap_bram_oarg_6_en0),
        .ap_bram_6_addr1(ap_bram_oarg_6_addr1),
        .ap_bram_6_din1(ap_bram_oarg_6_din1),
        .ap_bram_6_dout1(ap_bram_oarg_6_dout1),
        .ap_bram_6_we1(ap_bram_oarg_6_we1),
        .ap_bram_6_en1(ap_bram_oarg_6_en1),
        .m_axis_bram_7_tlast(m_axis_bram_7_tlast),
        .m_axis_bram_7_tvalid(m_axis_bram_7_tvalid),
        .m_axis_bram_7_tkeep(m_axis_bram_7_tkeep),
        .m_axis_bram_7_tstrb(m_axis_bram_7_tstrb),
        .m_axis_bram_7_tdata(m_axis_bram_7_tdata),
        .m_axis_bram_7_tready(m_axis_bram_7_tready),
        .ap_bram_7_addr0(ap_bram_oarg_7_addr0),
        .ap_bram_7_din0(ap_bram_oarg_7_din0),
        .ap_bram_7_dout0(ap_bram_oarg_7_dout0),
        .ap_bram_7_we0(ap_bram_oarg_7_we0),
        .ap_bram_7_en0(ap_bram_oarg_7_en0),
        .ap_bram_7_addr1(ap_bram_oarg_7_addr1),
        .ap_bram_7_din1(ap_bram_oarg_7_din1),
        .ap_bram_7_dout1(ap_bram_oarg_7_dout1),
        .ap_bram_7_we1(ap_bram_oarg_7_we1),
        .ap_bram_7_en1(ap_bram_oarg_7_en1),
        .m_axis_bram_8_tlast(m_axis_bram_8_tlast),
        .m_axis_bram_8_tvalid(m_axis_bram_8_tvalid),
        .m_axis_bram_8_tkeep(m_axis_bram_8_tkeep),
        .m_axis_bram_8_tstrb(m_axis_bram_8_tstrb),
        .m_axis_bram_8_tdata(m_axis_bram_8_tdata),
        .m_axis_bram_8_tready(m_axis_bram_8_tready),
        .ap_bram_8_addr0(ap_bram_oarg_8_addr0),
        .ap_bram_8_din0(ap_bram_oarg_8_din0),
        .ap_bram_8_dout0(ap_bram_oarg_8_dout0),
        .ap_bram_8_we0(ap_bram_oarg_8_we0),
        .ap_bram_8_en0(ap_bram_oarg_8_en0),
        .ap_bram_8_addr1(ap_bram_oarg_8_addr1),
        .ap_bram_8_din1(ap_bram_oarg_8_din1),
        .ap_bram_8_dout1(ap_bram_oarg_8_dout1),
        .ap_bram_8_we1(ap_bram_oarg_8_we1),
        .ap_bram_8_en1(ap_bram_oarg_8_en1),
        .m_axis_bram_9_tlast(m_axis_bram_9_tlast),
        .m_axis_bram_9_tvalid(m_axis_bram_9_tvalid),
        .m_axis_bram_9_tkeep(m_axis_bram_9_tkeep),
        .m_axis_bram_9_tstrb(m_axis_bram_9_tstrb),
        .m_axis_bram_9_tdata(m_axis_bram_9_tdata),
        .m_axis_bram_9_tready(m_axis_bram_9_tready),
        .ap_bram_9_addr0(ap_bram_oarg_9_addr0),
        .ap_bram_9_din0(ap_bram_oarg_9_din0),
        .ap_bram_9_dout0(ap_bram_oarg_9_dout0),
        .ap_bram_9_we0(ap_bram_oarg_9_we0),
        .ap_bram_9_en0(ap_bram_oarg_9_en0),
        .ap_bram_9_addr1(ap_bram_oarg_9_addr1),
        .ap_bram_9_din1(ap_bram_oarg_9_din1),
        .ap_bram_9_dout1(ap_bram_oarg_9_dout1),
        .ap_bram_9_we1(ap_bram_oarg_9_we1),
        .ap_bram_9_en1(ap_bram_oarg_9_en1),
        .m_axis_bram_10_tlast(m_axis_bram_10_tlast),
        .m_axis_bram_10_tvalid(m_axis_bram_10_tvalid),
        .m_axis_bram_10_tkeep(m_axis_bram_10_tkeep),
        .m_axis_bram_10_tstrb(m_axis_bram_10_tstrb),
        .m_axis_bram_10_tdata(m_axis_bram_10_tdata),
        .m_axis_bram_10_tready(m_axis_bram_10_tready),
        .ap_bram_10_addr0(ap_bram_oarg_10_addr0),
        .ap_bram_10_din0(ap_bram_oarg_10_din0),
        .ap_bram_10_dout0(ap_bram_oarg_10_dout0),
        .ap_bram_10_we0(ap_bram_oarg_10_we0),
        .ap_bram_10_en0(ap_bram_oarg_10_en0),
        .ap_bram_10_addr1(ap_bram_oarg_10_addr1),
        .ap_bram_10_din1(ap_bram_oarg_10_din1),
        .ap_bram_10_dout1(ap_bram_oarg_10_dout1),
        .ap_bram_10_we1(ap_bram_oarg_10_we1),
        .ap_bram_10_en1(ap_bram_oarg_10_en1),
        .m_axis_bram_11_tlast(m_axis_bram_11_tlast),
        .m_axis_bram_11_tvalid(m_axis_bram_11_tvalid),
        .m_axis_bram_11_tkeep(m_axis_bram_11_tkeep),
        .m_axis_bram_11_tstrb(m_axis_bram_11_tstrb),
        .m_axis_bram_11_tdata(m_axis_bram_11_tdata),
        .m_axis_bram_11_tready(m_axis_bram_11_tready),
        .ap_bram_11_addr0(ap_bram_oarg_11_addr0),
        .ap_bram_11_din0(ap_bram_oarg_11_din0),
        .ap_bram_11_dout0(ap_bram_oarg_11_dout0),
        .ap_bram_11_we0(ap_bram_oarg_11_we0),
        .ap_bram_11_en0(ap_bram_oarg_11_en0),
        .ap_bram_11_addr1(ap_bram_oarg_11_addr1),
        .ap_bram_11_din1(ap_bram_oarg_11_din1),
        .ap_bram_11_dout1(ap_bram_oarg_11_dout1),
        .ap_bram_11_we1(ap_bram_oarg_11_we1),
        .ap_bram_11_en1(ap_bram_oarg_11_en1),
        .m_axis_bram_12_tlast(m_axis_bram_12_tlast),
        .m_axis_bram_12_tvalid(m_axis_bram_12_tvalid),
        .m_axis_bram_12_tkeep(m_axis_bram_12_tkeep),
        .m_axis_bram_12_tstrb(m_axis_bram_12_tstrb),
        .m_axis_bram_12_tdata(m_axis_bram_12_tdata),
        .m_axis_bram_12_tready(m_axis_bram_12_tready),
        .ap_bram_12_addr0(ap_bram_oarg_12_addr0),
        .ap_bram_12_din0(ap_bram_oarg_12_din0),
        .ap_bram_12_dout0(ap_bram_oarg_12_dout0),
        .ap_bram_12_we0(ap_bram_oarg_12_we0),
        .ap_bram_12_en0(ap_bram_oarg_12_en0),
        .ap_bram_12_addr1(ap_bram_oarg_12_addr1),
        .ap_bram_12_din1(ap_bram_oarg_12_din1),
        .ap_bram_12_dout1(ap_bram_oarg_12_dout1),
        .ap_bram_12_we1(ap_bram_oarg_12_we1),
        .ap_bram_12_en1(ap_bram_oarg_12_en1),
        .m_axis_bram_13_tlast(m_axis_bram_13_tlast),
        .m_axis_bram_13_tvalid(m_axis_bram_13_tvalid),
        .m_axis_bram_13_tkeep(m_axis_bram_13_tkeep),
        .m_axis_bram_13_tstrb(m_axis_bram_13_tstrb),
        .m_axis_bram_13_tdata(m_axis_bram_13_tdata),
        .m_axis_bram_13_tready(m_axis_bram_13_tready),
        .ap_bram_13_addr0(ap_bram_oarg_13_addr0),
        .ap_bram_13_din0(ap_bram_oarg_13_din0),
        .ap_bram_13_dout0(ap_bram_oarg_13_dout0),
        .ap_bram_13_we0(ap_bram_oarg_13_we0),
        .ap_bram_13_en0(ap_bram_oarg_13_en0),
        .ap_bram_13_addr1(ap_bram_oarg_13_addr1),
        .ap_bram_13_din1(ap_bram_oarg_13_din1),
        .ap_bram_13_dout1(ap_bram_oarg_13_dout1),
        .ap_bram_13_we1(ap_bram_oarg_13_we1),
        .ap_bram_13_en1(ap_bram_oarg_13_en1),
        .m_axis_bram_14_tlast(m_axis_bram_14_tlast),
        .m_axis_bram_14_tvalid(m_axis_bram_14_tvalid),
        .m_axis_bram_14_tkeep(m_axis_bram_14_tkeep),
        .m_axis_bram_14_tstrb(m_axis_bram_14_tstrb),
        .m_axis_bram_14_tdata(m_axis_bram_14_tdata),
        .m_axis_bram_14_tready(m_axis_bram_14_tready),
        .ap_bram_14_addr0(ap_bram_oarg_14_addr0),
        .ap_bram_14_din0(ap_bram_oarg_14_din0),
        .ap_bram_14_dout0(ap_bram_oarg_14_dout0),
        .ap_bram_14_we0(ap_bram_oarg_14_we0),
        .ap_bram_14_en0(ap_bram_oarg_14_en0),
        .ap_bram_14_addr1(ap_bram_oarg_14_addr1),
        .ap_bram_14_din1(ap_bram_oarg_14_din1),
        .ap_bram_14_dout1(ap_bram_oarg_14_dout1),
        .ap_bram_14_we1(ap_bram_oarg_14_we1),
        .ap_bram_14_en1(ap_bram_oarg_14_en1),
        .m_axis_bram_15_tlast(m_axis_bram_15_tlast),
        .m_axis_bram_15_tvalid(m_axis_bram_15_tvalid),
        .m_axis_bram_15_tkeep(m_axis_bram_15_tkeep),
        .m_axis_bram_15_tstrb(m_axis_bram_15_tstrb),
        .m_axis_bram_15_tdata(m_axis_bram_15_tdata),
        .m_axis_bram_15_tready(m_axis_bram_15_tready),
        .ap_bram_15_addr0(ap_bram_oarg_15_addr0),
        .ap_bram_15_din0(ap_bram_oarg_15_din0),
        .ap_bram_15_dout0(ap_bram_oarg_15_dout0),
        .ap_bram_15_we0(ap_bram_oarg_15_we0),
        .ap_bram_15_en0(ap_bram_oarg_15_en0),
        .ap_bram_15_addr1(ap_bram_oarg_15_addr1),
        .ap_bram_15_din1(ap_bram_oarg_15_din1),
        .ap_bram_15_dout1(ap_bram_oarg_15_dout1),
        .ap_bram_15_we1(ap_bram_oarg_15_we1),
        .ap_bram_15_en1(ap_bram_oarg_15_en1),
        .m_axis_bram_16_tlast(m_axis_bram_16_tlast),
        .m_axis_bram_16_tvalid(m_axis_bram_16_tvalid),
        .m_axis_bram_16_tkeep(m_axis_bram_16_tkeep),
        .m_axis_bram_16_tstrb(m_axis_bram_16_tstrb),
        .m_axis_bram_16_tdata(m_axis_bram_16_tdata),
        .m_axis_bram_16_tready(m_axis_bram_16_tready),
        .ap_bram_16_addr0(ap_bram_oarg_16_addr0),
        .ap_bram_16_din0(ap_bram_oarg_16_din0),
        .ap_bram_16_dout0(ap_bram_oarg_16_dout0),
        .ap_bram_16_we0(ap_bram_oarg_16_we0),
        .ap_bram_16_en0(ap_bram_oarg_16_en0),
        .ap_bram_16_addr1(ap_bram_oarg_16_addr1),
        .ap_bram_16_din1(ap_bram_oarg_16_din1),
        .ap_bram_16_dout1(ap_bram_oarg_16_dout1),
        .ap_bram_16_we1(ap_bram_oarg_16_we1),
        .ap_bram_16_en1(ap_bram_oarg_16_en1),
        .m_axis_bram_17_tlast(m_axis_bram_17_tlast),
        .m_axis_bram_17_tvalid(m_axis_bram_17_tvalid),
        .m_axis_bram_17_tkeep(m_axis_bram_17_tkeep),
        .m_axis_bram_17_tstrb(m_axis_bram_17_tstrb),
        .m_axis_bram_17_tdata(m_axis_bram_17_tdata),
        .m_axis_bram_17_tready(m_axis_bram_17_tready),
        .ap_bram_17_addr0(ap_bram_oarg_17_addr0),
        .ap_bram_17_din0(ap_bram_oarg_17_din0),
        .ap_bram_17_dout0(ap_bram_oarg_17_dout0),
        .ap_bram_17_we0(ap_bram_oarg_17_we0),
        .ap_bram_17_en0(ap_bram_oarg_17_en0),
        .ap_bram_17_addr1(ap_bram_oarg_17_addr1),
        .ap_bram_17_din1(ap_bram_oarg_17_din1),
        .ap_bram_17_dout1(ap_bram_oarg_17_dout1),
        .ap_bram_17_we1(ap_bram_oarg_17_we1),
        .ap_bram_17_en1(ap_bram_oarg_17_en1),
        .m_axis_bram_18_tlast(m_axis_bram_18_tlast),
        .m_axis_bram_18_tvalid(m_axis_bram_18_tvalid),
        .m_axis_bram_18_tkeep(m_axis_bram_18_tkeep),
        .m_axis_bram_18_tstrb(m_axis_bram_18_tstrb),
        .m_axis_bram_18_tdata(m_axis_bram_18_tdata),
        .m_axis_bram_18_tready(m_axis_bram_18_tready),
        .ap_bram_18_addr0(ap_bram_oarg_18_addr0),
        .ap_bram_18_din0(ap_bram_oarg_18_din0),
        .ap_bram_18_dout0(ap_bram_oarg_18_dout0),
        .ap_bram_18_we0(ap_bram_oarg_18_we0),
        .ap_bram_18_en0(ap_bram_oarg_18_en0),
        .ap_bram_18_addr1(ap_bram_oarg_18_addr1),
        .ap_bram_18_din1(ap_bram_oarg_18_din1),
        .ap_bram_18_dout1(ap_bram_oarg_18_dout1),
        .ap_bram_18_we1(ap_bram_oarg_18_we1),
        .ap_bram_18_en1(ap_bram_oarg_18_en1),
        .m_axis_bram_19_tlast(m_axis_bram_19_tlast),
        .m_axis_bram_19_tvalid(m_axis_bram_19_tvalid),
        .m_axis_bram_19_tkeep(m_axis_bram_19_tkeep),
        .m_axis_bram_19_tstrb(m_axis_bram_19_tstrb),
        .m_axis_bram_19_tdata(m_axis_bram_19_tdata),
        .m_axis_bram_19_tready(m_axis_bram_19_tready),
        .ap_bram_19_addr0(ap_bram_oarg_19_addr0),
        .ap_bram_19_din0(ap_bram_oarg_19_din0),
        .ap_bram_19_dout0(ap_bram_oarg_19_dout0),
        .ap_bram_19_we0(ap_bram_oarg_19_we0),
        .ap_bram_19_en0(ap_bram_oarg_19_en0),
        .ap_bram_19_addr1(ap_bram_oarg_19_addr1),
        .ap_bram_19_din1(ap_bram_oarg_19_din1),
        .ap_bram_19_dout1(ap_bram_oarg_19_dout1),
        .ap_bram_19_we1(ap_bram_oarg_19_we1),
        .ap_bram_19_en1(ap_bram_oarg_19_en1),
        .m_axis_bram_20_tlast(m_axis_bram_20_tlast),
        .m_axis_bram_20_tvalid(m_axis_bram_20_tvalid),
        .m_axis_bram_20_tkeep(m_axis_bram_20_tkeep),
        .m_axis_bram_20_tstrb(m_axis_bram_20_tstrb),
        .m_axis_bram_20_tdata(m_axis_bram_20_tdata),
        .m_axis_bram_20_tready(m_axis_bram_20_tready),
        .ap_bram_20_addr0(ap_bram_oarg_20_addr0),
        .ap_bram_20_din0(ap_bram_oarg_20_din0),
        .ap_bram_20_dout0(ap_bram_oarg_20_dout0),
        .ap_bram_20_we0(ap_bram_oarg_20_we0),
        .ap_bram_20_en0(ap_bram_oarg_20_en0),
        .ap_bram_20_addr1(ap_bram_oarg_20_addr1),
        .ap_bram_20_din1(ap_bram_oarg_20_din1),
        .ap_bram_20_dout1(ap_bram_oarg_20_dout1),
        .ap_bram_20_we1(ap_bram_oarg_20_we1),
        .ap_bram_20_en1(ap_bram_oarg_20_en1),
        .m_axis_bram_21_tlast(m_axis_bram_21_tlast),
        .m_axis_bram_21_tvalid(m_axis_bram_21_tvalid),
        .m_axis_bram_21_tkeep(m_axis_bram_21_tkeep),
        .m_axis_bram_21_tstrb(m_axis_bram_21_tstrb),
        .m_axis_bram_21_tdata(m_axis_bram_21_tdata),
        .m_axis_bram_21_tready(m_axis_bram_21_tready),
        .ap_bram_21_addr0(ap_bram_oarg_21_addr0),
        .ap_bram_21_din0(ap_bram_oarg_21_din0),
        .ap_bram_21_dout0(ap_bram_oarg_21_dout0),
        .ap_bram_21_we0(ap_bram_oarg_21_we0),
        .ap_bram_21_en0(ap_bram_oarg_21_en0),
        .ap_bram_21_addr1(ap_bram_oarg_21_addr1),
        .ap_bram_21_din1(ap_bram_oarg_21_din1),
        .ap_bram_21_dout1(ap_bram_oarg_21_dout1),
        .ap_bram_21_we1(ap_bram_oarg_21_we1),
        .ap_bram_21_en1(ap_bram_oarg_21_en1),
        .m_axis_bram_22_tlast(m_axis_bram_22_tlast),
        .m_axis_bram_22_tvalid(m_axis_bram_22_tvalid),
        .m_axis_bram_22_tkeep(m_axis_bram_22_tkeep),
        .m_axis_bram_22_tstrb(m_axis_bram_22_tstrb),
        .m_axis_bram_22_tdata(m_axis_bram_22_tdata),
        .m_axis_bram_22_tready(m_axis_bram_22_tready),
        .ap_bram_22_addr0(ap_bram_oarg_22_addr0),
        .ap_bram_22_din0(ap_bram_oarg_22_din0),
        .ap_bram_22_dout0(ap_bram_oarg_22_dout0),
        .ap_bram_22_we0(ap_bram_oarg_22_we0),
        .ap_bram_22_en0(ap_bram_oarg_22_en0),
        .ap_bram_22_addr1(ap_bram_oarg_22_addr1),
        .ap_bram_22_din1(ap_bram_oarg_22_din1),
        .ap_bram_22_dout1(ap_bram_oarg_22_dout1),
        .ap_bram_22_we1(ap_bram_oarg_22_we1),
        .ap_bram_22_en1(ap_bram_oarg_22_en1),
        .m_axis_bram_23_tlast(m_axis_bram_23_tlast),
        .m_axis_bram_23_tvalid(m_axis_bram_23_tvalid),
        .m_axis_bram_23_tkeep(m_axis_bram_23_tkeep),
        .m_axis_bram_23_tstrb(m_axis_bram_23_tstrb),
        .m_axis_bram_23_tdata(m_axis_bram_23_tdata),
        .m_axis_bram_23_tready(m_axis_bram_23_tready),
        .ap_bram_23_addr0(ap_bram_oarg_23_addr0),
        .ap_bram_23_din0(ap_bram_oarg_23_din0),
        .ap_bram_23_dout0(ap_bram_oarg_23_dout0),
        .ap_bram_23_we0(ap_bram_oarg_23_we0),
        .ap_bram_23_en0(ap_bram_oarg_23_en0),
        .ap_bram_23_addr1(ap_bram_oarg_23_addr1),
        .ap_bram_23_din1(ap_bram_oarg_23_din1),
        .ap_bram_23_dout1(ap_bram_oarg_23_dout1),
        .ap_bram_23_we1(ap_bram_oarg_23_we1),
        .ap_bram_23_en1(ap_bram_oarg_23_en1),
        .m_axis_bram_24_tlast(m_axis_bram_24_tlast),
        .m_axis_bram_24_tvalid(m_axis_bram_24_tvalid),
        .m_axis_bram_24_tkeep(m_axis_bram_24_tkeep),
        .m_axis_bram_24_tstrb(m_axis_bram_24_tstrb),
        .m_axis_bram_24_tdata(m_axis_bram_24_tdata),
        .m_axis_bram_24_tready(m_axis_bram_24_tready),
        .ap_bram_24_addr0(ap_bram_oarg_24_addr0),
        .ap_bram_24_din0(ap_bram_oarg_24_din0),
        .ap_bram_24_dout0(ap_bram_oarg_24_dout0),
        .ap_bram_24_we0(ap_bram_oarg_24_we0),
        .ap_bram_24_en0(ap_bram_oarg_24_en0),
        .ap_bram_24_addr1(ap_bram_oarg_24_addr1),
        .ap_bram_24_din1(ap_bram_oarg_24_din1),
        .ap_bram_24_dout1(ap_bram_oarg_24_dout1),
        .ap_bram_24_we1(ap_bram_oarg_24_we1),
        .ap_bram_24_en1(ap_bram_oarg_24_en1),
        .m_axis_bram_25_tlast(m_axis_bram_25_tlast),
        .m_axis_bram_25_tvalid(m_axis_bram_25_tvalid),
        .m_axis_bram_25_tkeep(m_axis_bram_25_tkeep),
        .m_axis_bram_25_tstrb(m_axis_bram_25_tstrb),
        .m_axis_bram_25_tdata(m_axis_bram_25_tdata),
        .m_axis_bram_25_tready(m_axis_bram_25_tready),
        .ap_bram_25_addr0(ap_bram_oarg_25_addr0),
        .ap_bram_25_din0(ap_bram_oarg_25_din0),
        .ap_bram_25_dout0(ap_bram_oarg_25_dout0),
        .ap_bram_25_we0(ap_bram_oarg_25_we0),
        .ap_bram_25_en0(ap_bram_oarg_25_en0),
        .ap_bram_25_addr1(ap_bram_oarg_25_addr1),
        .ap_bram_25_din1(ap_bram_oarg_25_din1),
        .ap_bram_25_dout1(ap_bram_oarg_25_dout1),
        .ap_bram_25_we1(ap_bram_oarg_25_we1),
        .ap_bram_25_en1(ap_bram_oarg_25_en1),
        .m_axis_bram_26_tlast(m_axis_bram_26_tlast),
        .m_axis_bram_26_tvalid(m_axis_bram_26_tvalid),
        .m_axis_bram_26_tkeep(m_axis_bram_26_tkeep),
        .m_axis_bram_26_tstrb(m_axis_bram_26_tstrb),
        .m_axis_bram_26_tdata(m_axis_bram_26_tdata),
        .m_axis_bram_26_tready(m_axis_bram_26_tready),
        .ap_bram_26_addr0(ap_bram_oarg_26_addr0),
        .ap_bram_26_din0(ap_bram_oarg_26_din0),
        .ap_bram_26_dout0(ap_bram_oarg_26_dout0),
        .ap_bram_26_we0(ap_bram_oarg_26_we0),
        .ap_bram_26_en0(ap_bram_oarg_26_en0),
        .ap_bram_26_addr1(ap_bram_oarg_26_addr1),
        .ap_bram_26_din1(ap_bram_oarg_26_din1),
        .ap_bram_26_dout1(ap_bram_oarg_26_dout1),
        .ap_bram_26_we1(ap_bram_oarg_26_we1),
        .ap_bram_26_en1(ap_bram_oarg_26_en1),
        .m_axis_bram_27_tlast(m_axis_bram_27_tlast),
        .m_axis_bram_27_tvalid(m_axis_bram_27_tvalid),
        .m_axis_bram_27_tkeep(m_axis_bram_27_tkeep),
        .m_axis_bram_27_tstrb(m_axis_bram_27_tstrb),
        .m_axis_bram_27_tdata(m_axis_bram_27_tdata),
        .m_axis_bram_27_tready(m_axis_bram_27_tready),
        .ap_bram_27_addr0(ap_bram_oarg_27_addr0),
        .ap_bram_27_din0(ap_bram_oarg_27_din0),
        .ap_bram_27_dout0(ap_bram_oarg_27_dout0),
        .ap_bram_27_we0(ap_bram_oarg_27_we0),
        .ap_bram_27_en0(ap_bram_oarg_27_en0),
        .ap_bram_27_addr1(ap_bram_oarg_27_addr1),
        .ap_bram_27_din1(ap_bram_oarg_27_din1),
        .ap_bram_27_dout1(ap_bram_oarg_27_dout1),
        .ap_bram_27_we1(ap_bram_oarg_27_we1),
        .ap_bram_27_en1(ap_bram_oarg_27_en1),
        .m_axis_bram_28_tlast(m_axis_bram_28_tlast),
        .m_axis_bram_28_tvalid(m_axis_bram_28_tvalid),
        .m_axis_bram_28_tkeep(m_axis_bram_28_tkeep),
        .m_axis_bram_28_tstrb(m_axis_bram_28_tstrb),
        .m_axis_bram_28_tdata(m_axis_bram_28_tdata),
        .m_axis_bram_28_tready(m_axis_bram_28_tready),
        .ap_bram_28_addr0(ap_bram_oarg_28_addr0),
        .ap_bram_28_din0(ap_bram_oarg_28_din0),
        .ap_bram_28_dout0(ap_bram_oarg_28_dout0),
        .ap_bram_28_we0(ap_bram_oarg_28_we0),
        .ap_bram_28_en0(ap_bram_oarg_28_en0),
        .ap_bram_28_addr1(ap_bram_oarg_28_addr1),
        .ap_bram_28_din1(ap_bram_oarg_28_din1),
        .ap_bram_28_dout1(ap_bram_oarg_28_dout1),
        .ap_bram_28_we1(ap_bram_oarg_28_we1),
        .ap_bram_28_en1(ap_bram_oarg_28_en1),
        .m_axis_bram_29_tlast(m_axis_bram_29_tlast),
        .m_axis_bram_29_tvalid(m_axis_bram_29_tvalid),
        .m_axis_bram_29_tkeep(m_axis_bram_29_tkeep),
        .m_axis_bram_29_tstrb(m_axis_bram_29_tstrb),
        .m_axis_bram_29_tdata(m_axis_bram_29_tdata),
        .m_axis_bram_29_tready(m_axis_bram_29_tready),
        .ap_bram_29_addr0(ap_bram_oarg_29_addr0),
        .ap_bram_29_din0(ap_bram_oarg_29_din0),
        .ap_bram_29_dout0(ap_bram_oarg_29_dout0),
        .ap_bram_29_we0(ap_bram_oarg_29_we0),
        .ap_bram_29_en0(ap_bram_oarg_29_en0),
        .ap_bram_29_addr1(ap_bram_oarg_29_addr1),
        .ap_bram_29_din1(ap_bram_oarg_29_din1),
        .ap_bram_29_dout1(ap_bram_oarg_29_dout1),
        .ap_bram_29_we1(ap_bram_oarg_29_we1),
        .ap_bram_29_en1(ap_bram_oarg_29_en1),
        .m_axis_bram_30_tlast(m_axis_bram_30_tlast),
        .m_axis_bram_30_tvalid(m_axis_bram_30_tvalid),
        .m_axis_bram_30_tkeep(m_axis_bram_30_tkeep),
        .m_axis_bram_30_tstrb(m_axis_bram_30_tstrb),
        .m_axis_bram_30_tdata(m_axis_bram_30_tdata),
        .m_axis_bram_30_tready(m_axis_bram_30_tready),
        .ap_bram_30_addr0(ap_bram_oarg_30_addr0),
        .ap_bram_30_din0(ap_bram_oarg_30_din0),
        .ap_bram_30_dout0(ap_bram_oarg_30_dout0),
        .ap_bram_30_we0(ap_bram_oarg_30_we0),
        .ap_bram_30_en0(ap_bram_oarg_30_en0),
        .ap_bram_30_addr1(ap_bram_oarg_30_addr1),
        .ap_bram_30_din1(ap_bram_oarg_30_din1),
        .ap_bram_30_dout1(ap_bram_oarg_30_dout1),
        .ap_bram_30_we1(ap_bram_oarg_30_we1),
        .ap_bram_30_en1(ap_bram_oarg_30_en1),
        .m_axis_bram_31_tlast(m_axis_bram_31_tlast),
        .m_axis_bram_31_tvalid(m_axis_bram_31_tvalid),
        .m_axis_bram_31_tkeep(m_axis_bram_31_tkeep),
        .m_axis_bram_31_tstrb(m_axis_bram_31_tstrb),
        .m_axis_bram_31_tdata(m_axis_bram_31_tdata),
        .m_axis_bram_31_tready(m_axis_bram_31_tready),
        .ap_bram_31_addr0(ap_bram_oarg_31_addr0),
        .ap_bram_31_din0(ap_bram_oarg_31_din0),
        .ap_bram_31_dout0(ap_bram_oarg_31_dout0),
        .ap_bram_31_we0(ap_bram_oarg_31_we0),
        .ap_bram_31_en0(ap_bram_oarg_31_en0),
        .ap_bram_31_addr1(ap_bram_oarg_31_addr1),
        .ap_bram_31_din1(ap_bram_oarg_31_din1),
        .ap_bram_31_dout1(ap_bram_oarg_31_dout1),
        .ap_bram_31_we1(ap_bram_oarg_31_we1),
        .ap_bram_31_en1(ap_bram_oarg_31_en1),
        .m_axis_bram_32_tlast(m_axis_bram_32_tlast),
        .m_axis_bram_32_tvalid(m_axis_bram_32_tvalid),
        .m_axis_bram_32_tkeep(m_axis_bram_32_tkeep),
        .m_axis_bram_32_tstrb(m_axis_bram_32_tstrb),
        .m_axis_bram_32_tdata(m_axis_bram_32_tdata),
        .m_axis_bram_32_tready(m_axis_bram_32_tready),
        .ap_bram_32_addr0(ap_bram_oarg_32_addr0),
        .ap_bram_32_din0(ap_bram_oarg_32_din0),
        .ap_bram_32_dout0(ap_bram_oarg_32_dout0),
        .ap_bram_32_we0(ap_bram_oarg_32_we0),
        .ap_bram_32_en0(ap_bram_oarg_32_en0),
        .ap_bram_32_addr1(ap_bram_oarg_32_addr1),
        .ap_bram_32_din1(ap_bram_oarg_32_din1),
        .ap_bram_32_dout1(ap_bram_oarg_32_dout1),
        .ap_bram_32_we1(ap_bram_oarg_32_we1),
        .ap_bram_32_en1(ap_bram_oarg_32_en1),
        .m_axis_bram_33_tlast(m_axis_bram_33_tlast),
        .m_axis_bram_33_tvalid(m_axis_bram_33_tvalid),
        .m_axis_bram_33_tkeep(m_axis_bram_33_tkeep),
        .m_axis_bram_33_tstrb(m_axis_bram_33_tstrb),
        .m_axis_bram_33_tdata(m_axis_bram_33_tdata),
        .m_axis_bram_33_tready(m_axis_bram_33_tready),
        .ap_bram_33_addr0(ap_bram_oarg_33_addr0),
        .ap_bram_33_din0(ap_bram_oarg_33_din0),
        .ap_bram_33_dout0(ap_bram_oarg_33_dout0),
        .ap_bram_33_we0(ap_bram_oarg_33_we0),
        .ap_bram_33_en0(ap_bram_oarg_33_en0),
        .ap_bram_33_addr1(ap_bram_oarg_33_addr1),
        .ap_bram_33_din1(ap_bram_oarg_33_din1),
        .ap_bram_33_dout1(ap_bram_oarg_33_dout1),
        .ap_bram_33_we1(ap_bram_oarg_33_we1),
        .ap_bram_33_en1(ap_bram_oarg_33_en1),
        .m_axis_bram_34_tlast(m_axis_bram_34_tlast),
        .m_axis_bram_34_tvalid(m_axis_bram_34_tvalid),
        .m_axis_bram_34_tkeep(m_axis_bram_34_tkeep),
        .m_axis_bram_34_tstrb(m_axis_bram_34_tstrb),
        .m_axis_bram_34_tdata(m_axis_bram_34_tdata),
        .m_axis_bram_34_tready(m_axis_bram_34_tready),
        .ap_bram_34_addr0(ap_bram_oarg_34_addr0),
        .ap_bram_34_din0(ap_bram_oarg_34_din0),
        .ap_bram_34_dout0(ap_bram_oarg_34_dout0),
        .ap_bram_34_we0(ap_bram_oarg_34_we0),
        .ap_bram_34_en0(ap_bram_oarg_34_en0),
        .ap_bram_34_addr1(ap_bram_oarg_34_addr1),
        .ap_bram_34_din1(ap_bram_oarg_34_din1),
        .ap_bram_34_dout1(ap_bram_oarg_34_dout1),
        .ap_bram_34_we1(ap_bram_oarg_34_we1),
        .ap_bram_34_en1(ap_bram_oarg_34_en1),
        .m_axis_bram_35_tlast(m_axis_bram_35_tlast),
        .m_axis_bram_35_tvalid(m_axis_bram_35_tvalid),
        .m_axis_bram_35_tkeep(m_axis_bram_35_tkeep),
        .m_axis_bram_35_tstrb(m_axis_bram_35_tstrb),
        .m_axis_bram_35_tdata(m_axis_bram_35_tdata),
        .m_axis_bram_35_tready(m_axis_bram_35_tready),
        .ap_bram_35_addr0(ap_bram_oarg_35_addr0),
        .ap_bram_35_din0(ap_bram_oarg_35_din0),
        .ap_bram_35_dout0(ap_bram_oarg_35_dout0),
        .ap_bram_35_we0(ap_bram_oarg_35_we0),
        .ap_bram_35_en0(ap_bram_oarg_35_en0),
        .ap_bram_35_addr1(ap_bram_oarg_35_addr1),
        .ap_bram_35_din1(ap_bram_oarg_35_din1),
        .ap_bram_35_dout1(ap_bram_oarg_35_dout1),
        .ap_bram_35_we1(ap_bram_oarg_35_we1),
        .ap_bram_35_en1(ap_bram_oarg_35_en1),
        .m_axis_bram_36_tlast(m_axis_bram_36_tlast),
        .m_axis_bram_36_tvalid(m_axis_bram_36_tvalid),
        .m_axis_bram_36_tkeep(m_axis_bram_36_tkeep),
        .m_axis_bram_36_tstrb(m_axis_bram_36_tstrb),
        .m_axis_bram_36_tdata(m_axis_bram_36_tdata),
        .m_axis_bram_36_tready(m_axis_bram_36_tready),
        .ap_bram_36_addr0(ap_bram_oarg_36_addr0),
        .ap_bram_36_din0(ap_bram_oarg_36_din0),
        .ap_bram_36_dout0(ap_bram_oarg_36_dout0),
        .ap_bram_36_we0(ap_bram_oarg_36_we0),
        .ap_bram_36_en0(ap_bram_oarg_36_en0),
        .ap_bram_36_addr1(ap_bram_oarg_36_addr1),
        .ap_bram_36_din1(ap_bram_oarg_36_din1),
        .ap_bram_36_dout1(ap_bram_oarg_36_dout1),
        .ap_bram_36_we1(ap_bram_oarg_36_we1),
        .ap_bram_36_en1(ap_bram_oarg_36_en1),
        .m_axis_bram_37_tlast(m_axis_bram_37_tlast),
        .m_axis_bram_37_tvalid(m_axis_bram_37_tvalid),
        .m_axis_bram_37_tkeep(m_axis_bram_37_tkeep),
        .m_axis_bram_37_tstrb(m_axis_bram_37_tstrb),
        .m_axis_bram_37_tdata(m_axis_bram_37_tdata),
        .m_axis_bram_37_tready(m_axis_bram_37_tready),
        .ap_bram_37_addr0(ap_bram_oarg_37_addr0),
        .ap_bram_37_din0(ap_bram_oarg_37_din0),
        .ap_bram_37_dout0(ap_bram_oarg_37_dout0),
        .ap_bram_37_we0(ap_bram_oarg_37_we0),
        .ap_bram_37_en0(ap_bram_oarg_37_en0),
        .ap_bram_37_addr1(ap_bram_oarg_37_addr1),
        .ap_bram_37_din1(ap_bram_oarg_37_din1),
        .ap_bram_37_dout1(ap_bram_oarg_37_dout1),
        .ap_bram_37_we1(ap_bram_oarg_37_we1),
        .ap_bram_37_en1(ap_bram_oarg_37_en1),
        .m_axis_bram_38_tlast(m_axis_bram_38_tlast),
        .m_axis_bram_38_tvalid(m_axis_bram_38_tvalid),
        .m_axis_bram_38_tkeep(m_axis_bram_38_tkeep),
        .m_axis_bram_38_tstrb(m_axis_bram_38_tstrb),
        .m_axis_bram_38_tdata(m_axis_bram_38_tdata),
        .m_axis_bram_38_tready(m_axis_bram_38_tready),
        .ap_bram_38_addr0(ap_bram_oarg_38_addr0),
        .ap_bram_38_din0(ap_bram_oarg_38_din0),
        .ap_bram_38_dout0(ap_bram_oarg_38_dout0),
        .ap_bram_38_we0(ap_bram_oarg_38_we0),
        .ap_bram_38_en0(ap_bram_oarg_38_en0),
        .ap_bram_38_addr1(ap_bram_oarg_38_addr1),
        .ap_bram_38_din1(ap_bram_oarg_38_din1),
        .ap_bram_38_dout1(ap_bram_oarg_38_dout1),
        .ap_bram_38_we1(ap_bram_oarg_38_we1),
        .ap_bram_38_en1(ap_bram_oarg_38_en1),
        .m_axis_bram_39_tlast(m_axis_bram_39_tlast),
        .m_axis_bram_39_tvalid(m_axis_bram_39_tvalid),
        .m_axis_bram_39_tkeep(m_axis_bram_39_tkeep),
        .m_axis_bram_39_tstrb(m_axis_bram_39_tstrb),
        .m_axis_bram_39_tdata(m_axis_bram_39_tdata),
        .m_axis_bram_39_tready(m_axis_bram_39_tready),
        .ap_bram_39_addr0(ap_bram_oarg_39_addr0),
        .ap_bram_39_din0(ap_bram_oarg_39_din0),
        .ap_bram_39_dout0(ap_bram_oarg_39_dout0),
        .ap_bram_39_we0(ap_bram_oarg_39_we0),
        .ap_bram_39_en0(ap_bram_oarg_39_en0),
        .ap_bram_39_addr1(ap_bram_oarg_39_addr1),
        .ap_bram_39_din1(ap_bram_oarg_39_din1),
        .ap_bram_39_dout1(ap_bram_oarg_39_dout1),
        .ap_bram_39_we1(ap_bram_oarg_39_we1),
        .ap_bram_39_en1(ap_bram_oarg_39_en1),
        .m_axis_bram_40_tlast(m_axis_bram_40_tlast),
        .m_axis_bram_40_tvalid(m_axis_bram_40_tvalid),
        .m_axis_bram_40_tkeep(m_axis_bram_40_tkeep),
        .m_axis_bram_40_tstrb(m_axis_bram_40_tstrb),
        .m_axis_bram_40_tdata(m_axis_bram_40_tdata),
        .m_axis_bram_40_tready(m_axis_bram_40_tready),
        .ap_bram_40_addr0(ap_bram_oarg_40_addr0),
        .ap_bram_40_din0(ap_bram_oarg_40_din0),
        .ap_bram_40_dout0(ap_bram_oarg_40_dout0),
        .ap_bram_40_we0(ap_bram_oarg_40_we0),
        .ap_bram_40_en0(ap_bram_oarg_40_en0),
        .ap_bram_40_addr1(ap_bram_oarg_40_addr1),
        .ap_bram_40_din1(ap_bram_oarg_40_din1),
        .ap_bram_40_dout1(ap_bram_oarg_40_dout1),
        .ap_bram_40_we1(ap_bram_oarg_40_we1),
        .ap_bram_40_en1(ap_bram_oarg_40_en1),
        .m_axis_bram_41_tlast(m_axis_bram_41_tlast),
        .m_axis_bram_41_tvalid(m_axis_bram_41_tvalid),
        .m_axis_bram_41_tkeep(m_axis_bram_41_tkeep),
        .m_axis_bram_41_tstrb(m_axis_bram_41_tstrb),
        .m_axis_bram_41_tdata(m_axis_bram_41_tdata),
        .m_axis_bram_41_tready(m_axis_bram_41_tready),
        .ap_bram_41_addr0(ap_bram_oarg_41_addr0),
        .ap_bram_41_din0(ap_bram_oarg_41_din0),
        .ap_bram_41_dout0(ap_bram_oarg_41_dout0),
        .ap_bram_41_we0(ap_bram_oarg_41_we0),
        .ap_bram_41_en0(ap_bram_oarg_41_en0),
        .ap_bram_41_addr1(ap_bram_oarg_41_addr1),
        .ap_bram_41_din1(ap_bram_oarg_41_din1),
        .ap_bram_41_dout1(ap_bram_oarg_41_dout1),
        .ap_bram_41_we1(ap_bram_oarg_41_we1),
        .ap_bram_41_en1(ap_bram_oarg_41_en1),
        .m_axis_bram_42_tlast(m_axis_bram_42_tlast),
        .m_axis_bram_42_tvalid(m_axis_bram_42_tvalid),
        .m_axis_bram_42_tkeep(m_axis_bram_42_tkeep),
        .m_axis_bram_42_tstrb(m_axis_bram_42_tstrb),
        .m_axis_bram_42_tdata(m_axis_bram_42_tdata),
        .m_axis_bram_42_tready(m_axis_bram_42_tready),
        .ap_bram_42_addr0(ap_bram_oarg_42_addr0),
        .ap_bram_42_din0(ap_bram_oarg_42_din0),
        .ap_bram_42_dout0(ap_bram_oarg_42_dout0),
        .ap_bram_42_we0(ap_bram_oarg_42_we0),
        .ap_bram_42_en0(ap_bram_oarg_42_en0),
        .ap_bram_42_addr1(ap_bram_oarg_42_addr1),
        .ap_bram_42_din1(ap_bram_oarg_42_din1),
        .ap_bram_42_dout1(ap_bram_oarg_42_dout1),
        .ap_bram_42_we1(ap_bram_oarg_42_we1),
        .ap_bram_42_en1(ap_bram_oarg_42_en1),
        .m_axis_bram_43_tlast(m_axis_bram_43_tlast),
        .m_axis_bram_43_tvalid(m_axis_bram_43_tvalid),
        .m_axis_bram_43_tkeep(m_axis_bram_43_tkeep),
        .m_axis_bram_43_tstrb(m_axis_bram_43_tstrb),
        .m_axis_bram_43_tdata(m_axis_bram_43_tdata),
        .m_axis_bram_43_tready(m_axis_bram_43_tready),
        .ap_bram_43_addr0(ap_bram_oarg_43_addr0),
        .ap_bram_43_din0(ap_bram_oarg_43_din0),
        .ap_bram_43_dout0(ap_bram_oarg_43_dout0),
        .ap_bram_43_we0(ap_bram_oarg_43_we0),
        .ap_bram_43_en0(ap_bram_oarg_43_en0),
        .ap_bram_43_addr1(ap_bram_oarg_43_addr1),
        .ap_bram_43_din1(ap_bram_oarg_43_din1),
        .ap_bram_43_dout1(ap_bram_oarg_43_dout1),
        .ap_bram_43_we1(ap_bram_oarg_43_we1),
        .ap_bram_43_en1(ap_bram_oarg_43_en1),
        .m_axis_bram_44_tlast(m_axis_bram_44_tlast),
        .m_axis_bram_44_tvalid(m_axis_bram_44_tvalid),
        .m_axis_bram_44_tkeep(m_axis_bram_44_tkeep),
        .m_axis_bram_44_tstrb(m_axis_bram_44_tstrb),
        .m_axis_bram_44_tdata(m_axis_bram_44_tdata),
        .m_axis_bram_44_tready(m_axis_bram_44_tready),
        .ap_bram_44_addr0(ap_bram_oarg_44_addr0),
        .ap_bram_44_din0(ap_bram_oarg_44_din0),
        .ap_bram_44_dout0(ap_bram_oarg_44_dout0),
        .ap_bram_44_we0(ap_bram_oarg_44_we0),
        .ap_bram_44_en0(ap_bram_oarg_44_en0),
        .ap_bram_44_addr1(ap_bram_oarg_44_addr1),
        .ap_bram_44_din1(ap_bram_oarg_44_din1),
        .ap_bram_44_dout1(ap_bram_oarg_44_dout1),
        .ap_bram_44_we1(ap_bram_oarg_44_we1),
        .ap_bram_44_en1(ap_bram_oarg_44_en1),
        .m_axis_bram_45_tlast(m_axis_bram_45_tlast),
        .m_axis_bram_45_tvalid(m_axis_bram_45_tvalid),
        .m_axis_bram_45_tkeep(m_axis_bram_45_tkeep),
        .m_axis_bram_45_tstrb(m_axis_bram_45_tstrb),
        .m_axis_bram_45_tdata(m_axis_bram_45_tdata),
        .m_axis_bram_45_tready(m_axis_bram_45_tready),
        .ap_bram_45_addr0(ap_bram_oarg_45_addr0),
        .ap_bram_45_din0(ap_bram_oarg_45_din0),
        .ap_bram_45_dout0(ap_bram_oarg_45_dout0),
        .ap_bram_45_we0(ap_bram_oarg_45_we0),
        .ap_bram_45_en0(ap_bram_oarg_45_en0),
        .ap_bram_45_addr1(ap_bram_oarg_45_addr1),
        .ap_bram_45_din1(ap_bram_oarg_45_din1),
        .ap_bram_45_dout1(ap_bram_oarg_45_dout1),
        .ap_bram_45_we1(ap_bram_oarg_45_we1),
        .ap_bram_45_en1(ap_bram_oarg_45_en1),
        .m_axis_bram_46_tlast(m_axis_bram_46_tlast),
        .m_axis_bram_46_tvalid(m_axis_bram_46_tvalid),
        .m_axis_bram_46_tkeep(m_axis_bram_46_tkeep),
        .m_axis_bram_46_tstrb(m_axis_bram_46_tstrb),
        .m_axis_bram_46_tdata(m_axis_bram_46_tdata),
        .m_axis_bram_46_tready(m_axis_bram_46_tready),
        .ap_bram_46_addr0(ap_bram_oarg_46_addr0),
        .ap_bram_46_din0(ap_bram_oarg_46_din0),
        .ap_bram_46_dout0(ap_bram_oarg_46_dout0),
        .ap_bram_46_we0(ap_bram_oarg_46_we0),
        .ap_bram_46_en0(ap_bram_oarg_46_en0),
        .ap_bram_46_addr1(ap_bram_oarg_46_addr1),
        .ap_bram_46_din1(ap_bram_oarg_46_din1),
        .ap_bram_46_dout1(ap_bram_oarg_46_dout1),
        .ap_bram_46_we1(ap_bram_oarg_46_we1),
        .ap_bram_46_en1(ap_bram_oarg_46_en1),
        .m_axis_bram_47_tlast(m_axis_bram_47_tlast),
        .m_axis_bram_47_tvalid(m_axis_bram_47_tvalid),
        .m_axis_bram_47_tkeep(m_axis_bram_47_tkeep),
        .m_axis_bram_47_tstrb(m_axis_bram_47_tstrb),
        .m_axis_bram_47_tdata(m_axis_bram_47_tdata),
        .m_axis_bram_47_tready(m_axis_bram_47_tready),
        .ap_bram_47_addr0(ap_bram_oarg_47_addr0),
        .ap_bram_47_din0(ap_bram_oarg_47_din0),
        .ap_bram_47_dout0(ap_bram_oarg_47_dout0),
        .ap_bram_47_we0(ap_bram_oarg_47_we0),
        .ap_bram_47_en0(ap_bram_oarg_47_en0),
        .ap_bram_47_addr1(ap_bram_oarg_47_addr1),
        .ap_bram_47_din1(ap_bram_oarg_47_din1),
        .ap_bram_47_dout1(ap_bram_oarg_47_dout1),
        .ap_bram_47_we1(ap_bram_oarg_47_we1),
        .ap_bram_47_en1(ap_bram_oarg_47_en1),
        .m_axis_bram_48_tlast(m_axis_bram_48_tlast),
        .m_axis_bram_48_tvalid(m_axis_bram_48_tvalid),
        .m_axis_bram_48_tkeep(m_axis_bram_48_tkeep),
        .m_axis_bram_48_tstrb(m_axis_bram_48_tstrb),
        .m_axis_bram_48_tdata(m_axis_bram_48_tdata),
        .m_axis_bram_48_tready(m_axis_bram_48_tready),
        .ap_bram_48_addr0(ap_bram_oarg_48_addr0),
        .ap_bram_48_din0(ap_bram_oarg_48_din0),
        .ap_bram_48_dout0(ap_bram_oarg_48_dout0),
        .ap_bram_48_we0(ap_bram_oarg_48_we0),
        .ap_bram_48_en0(ap_bram_oarg_48_en0),
        .ap_bram_48_addr1(ap_bram_oarg_48_addr1),
        .ap_bram_48_din1(ap_bram_oarg_48_din1),
        .ap_bram_48_dout1(ap_bram_oarg_48_dout1),
        .ap_bram_48_we1(ap_bram_oarg_48_we1),
        .ap_bram_48_en1(ap_bram_oarg_48_en1),
        .m_axis_bram_49_tlast(m_axis_bram_49_tlast),
        .m_axis_bram_49_tvalid(m_axis_bram_49_tvalid),
        .m_axis_bram_49_tkeep(m_axis_bram_49_tkeep),
        .m_axis_bram_49_tstrb(m_axis_bram_49_tstrb),
        .m_axis_bram_49_tdata(m_axis_bram_49_tdata),
        .m_axis_bram_49_tready(m_axis_bram_49_tready),
        .ap_bram_49_addr0(ap_bram_oarg_49_addr0),
        .ap_bram_49_din0(ap_bram_oarg_49_din0),
        .ap_bram_49_dout0(ap_bram_oarg_49_dout0),
        .ap_bram_49_we0(ap_bram_oarg_49_we0),
        .ap_bram_49_en0(ap_bram_oarg_49_en0),
        .ap_bram_49_addr1(ap_bram_oarg_49_addr1),
        .ap_bram_49_din1(ap_bram_oarg_49_din1),
        .ap_bram_49_dout1(ap_bram_oarg_49_dout1),
        .ap_bram_49_we1(ap_bram_oarg_49_we1),
        .ap_bram_49_en1(ap_bram_oarg_49_en1),
        .m_axis_bram_50_tlast(m_axis_bram_50_tlast),
        .m_axis_bram_50_tvalid(m_axis_bram_50_tvalid),
        .m_axis_bram_50_tkeep(m_axis_bram_50_tkeep),
        .m_axis_bram_50_tstrb(m_axis_bram_50_tstrb),
        .m_axis_bram_50_tdata(m_axis_bram_50_tdata),
        .m_axis_bram_50_tready(m_axis_bram_50_tready),
        .ap_bram_50_addr0(ap_bram_oarg_50_addr0),
        .ap_bram_50_din0(ap_bram_oarg_50_din0),
        .ap_bram_50_dout0(ap_bram_oarg_50_dout0),
        .ap_bram_50_we0(ap_bram_oarg_50_we0),
        .ap_bram_50_en0(ap_bram_oarg_50_en0),
        .ap_bram_50_addr1(ap_bram_oarg_50_addr1),
        .ap_bram_50_din1(ap_bram_oarg_50_din1),
        .ap_bram_50_dout1(ap_bram_oarg_50_dout1),
        .ap_bram_50_we1(ap_bram_oarg_50_we1),
        .ap_bram_50_en1(ap_bram_oarg_50_en1),
        .m_axis_bram_51_tlast(m_axis_bram_51_tlast),
        .m_axis_bram_51_tvalid(m_axis_bram_51_tvalid),
        .m_axis_bram_51_tkeep(m_axis_bram_51_tkeep),
        .m_axis_bram_51_tstrb(m_axis_bram_51_tstrb),
        .m_axis_bram_51_tdata(m_axis_bram_51_tdata),
        .m_axis_bram_51_tready(m_axis_bram_51_tready),
        .ap_bram_51_addr0(ap_bram_oarg_51_addr0),
        .ap_bram_51_din0(ap_bram_oarg_51_din0),
        .ap_bram_51_dout0(ap_bram_oarg_51_dout0),
        .ap_bram_51_we0(ap_bram_oarg_51_we0),
        .ap_bram_51_en0(ap_bram_oarg_51_en0),
        .ap_bram_51_addr1(ap_bram_oarg_51_addr1),
        .ap_bram_51_din1(ap_bram_oarg_51_din1),
        .ap_bram_51_dout1(ap_bram_oarg_51_dout1),
        .ap_bram_51_we1(ap_bram_oarg_51_we1),
        .ap_bram_51_en1(ap_bram_oarg_51_en1),
        .m_axis_bram_52_tlast(m_axis_bram_52_tlast),
        .m_axis_bram_52_tvalid(m_axis_bram_52_tvalid),
        .m_axis_bram_52_tkeep(m_axis_bram_52_tkeep),
        .m_axis_bram_52_tstrb(m_axis_bram_52_tstrb),
        .m_axis_bram_52_tdata(m_axis_bram_52_tdata),
        .m_axis_bram_52_tready(m_axis_bram_52_tready),
        .ap_bram_52_addr0(ap_bram_oarg_52_addr0),
        .ap_bram_52_din0(ap_bram_oarg_52_din0),
        .ap_bram_52_dout0(ap_bram_oarg_52_dout0),
        .ap_bram_52_we0(ap_bram_oarg_52_we0),
        .ap_bram_52_en0(ap_bram_oarg_52_en0),
        .ap_bram_52_addr1(ap_bram_oarg_52_addr1),
        .ap_bram_52_din1(ap_bram_oarg_52_din1),
        .ap_bram_52_dout1(ap_bram_oarg_52_dout1),
        .ap_bram_52_we1(ap_bram_oarg_52_we1),
        .ap_bram_52_en1(ap_bram_oarg_52_en1),
        .m_axis_bram_53_tlast(m_axis_bram_53_tlast),
        .m_axis_bram_53_tvalid(m_axis_bram_53_tvalid),
        .m_axis_bram_53_tkeep(m_axis_bram_53_tkeep),
        .m_axis_bram_53_tstrb(m_axis_bram_53_tstrb),
        .m_axis_bram_53_tdata(m_axis_bram_53_tdata),
        .m_axis_bram_53_tready(m_axis_bram_53_tready),
        .ap_bram_53_addr0(ap_bram_oarg_53_addr0),
        .ap_bram_53_din0(ap_bram_oarg_53_din0),
        .ap_bram_53_dout0(ap_bram_oarg_53_dout0),
        .ap_bram_53_we0(ap_bram_oarg_53_we0),
        .ap_bram_53_en0(ap_bram_oarg_53_en0),
        .ap_bram_53_addr1(ap_bram_oarg_53_addr1),
        .ap_bram_53_din1(ap_bram_oarg_53_din1),
        .ap_bram_53_dout1(ap_bram_oarg_53_dout1),
        .ap_bram_53_we1(ap_bram_oarg_53_we1),
        .ap_bram_53_en1(ap_bram_oarg_53_en1),
        .m_axis_bram_54_tlast(m_axis_bram_54_tlast),
        .m_axis_bram_54_tvalid(m_axis_bram_54_tvalid),
        .m_axis_bram_54_tkeep(m_axis_bram_54_tkeep),
        .m_axis_bram_54_tstrb(m_axis_bram_54_tstrb),
        .m_axis_bram_54_tdata(m_axis_bram_54_tdata),
        .m_axis_bram_54_tready(m_axis_bram_54_tready),
        .ap_bram_54_addr0(ap_bram_oarg_54_addr0),
        .ap_bram_54_din0(ap_bram_oarg_54_din0),
        .ap_bram_54_dout0(ap_bram_oarg_54_dout0),
        .ap_bram_54_we0(ap_bram_oarg_54_we0),
        .ap_bram_54_en0(ap_bram_oarg_54_en0),
        .ap_bram_54_addr1(ap_bram_oarg_54_addr1),
        .ap_bram_54_din1(ap_bram_oarg_54_din1),
        .ap_bram_54_dout1(ap_bram_oarg_54_dout1),
        .ap_bram_54_we1(ap_bram_oarg_54_we1),
        .ap_bram_54_en1(ap_bram_oarg_54_en1),
        .m_axis_bram_55_tlast(m_axis_bram_55_tlast),
        .m_axis_bram_55_tvalid(m_axis_bram_55_tvalid),
        .m_axis_bram_55_tkeep(m_axis_bram_55_tkeep),
        .m_axis_bram_55_tstrb(m_axis_bram_55_tstrb),
        .m_axis_bram_55_tdata(m_axis_bram_55_tdata),
        .m_axis_bram_55_tready(m_axis_bram_55_tready),
        .ap_bram_55_addr0(ap_bram_oarg_55_addr0),
        .ap_bram_55_din0(ap_bram_oarg_55_din0),
        .ap_bram_55_dout0(ap_bram_oarg_55_dout0),
        .ap_bram_55_we0(ap_bram_oarg_55_we0),
        .ap_bram_55_en0(ap_bram_oarg_55_en0),
        .ap_bram_55_addr1(ap_bram_oarg_55_addr1),
        .ap_bram_55_din1(ap_bram_oarg_55_din1),
        .ap_bram_55_dout1(ap_bram_oarg_55_dout1),
        .ap_bram_55_we1(ap_bram_oarg_55_we1),
        .ap_bram_55_en1(ap_bram_oarg_55_en1),
        .m_axis_bram_56_tlast(m_axis_bram_56_tlast),
        .m_axis_bram_56_tvalid(m_axis_bram_56_tvalid),
        .m_axis_bram_56_tkeep(m_axis_bram_56_tkeep),
        .m_axis_bram_56_tstrb(m_axis_bram_56_tstrb),
        .m_axis_bram_56_tdata(m_axis_bram_56_tdata),
        .m_axis_bram_56_tready(m_axis_bram_56_tready),
        .ap_bram_56_addr0(ap_bram_oarg_56_addr0),
        .ap_bram_56_din0(ap_bram_oarg_56_din0),
        .ap_bram_56_dout0(ap_bram_oarg_56_dout0),
        .ap_bram_56_we0(ap_bram_oarg_56_we0),
        .ap_bram_56_en0(ap_bram_oarg_56_en0),
        .ap_bram_56_addr1(ap_bram_oarg_56_addr1),
        .ap_bram_56_din1(ap_bram_oarg_56_din1),
        .ap_bram_56_dout1(ap_bram_oarg_56_dout1),
        .ap_bram_56_we1(ap_bram_oarg_56_we1),
        .ap_bram_56_en1(ap_bram_oarg_56_en1),
        .m_axis_bram_57_tlast(m_axis_bram_57_tlast),
        .m_axis_bram_57_tvalid(m_axis_bram_57_tvalid),
        .m_axis_bram_57_tkeep(m_axis_bram_57_tkeep),
        .m_axis_bram_57_tstrb(m_axis_bram_57_tstrb),
        .m_axis_bram_57_tdata(m_axis_bram_57_tdata),
        .m_axis_bram_57_tready(m_axis_bram_57_tready),
        .ap_bram_57_addr0(ap_bram_oarg_57_addr0),
        .ap_bram_57_din0(ap_bram_oarg_57_din0),
        .ap_bram_57_dout0(ap_bram_oarg_57_dout0),
        .ap_bram_57_we0(ap_bram_oarg_57_we0),
        .ap_bram_57_en0(ap_bram_oarg_57_en0),
        .ap_bram_57_addr1(ap_bram_oarg_57_addr1),
        .ap_bram_57_din1(ap_bram_oarg_57_din1),
        .ap_bram_57_dout1(ap_bram_oarg_57_dout1),
        .ap_bram_57_we1(ap_bram_oarg_57_we1),
        .ap_bram_57_en1(ap_bram_oarg_57_en1),
        .m_axis_bram_58_tlast(m_axis_bram_58_tlast),
        .m_axis_bram_58_tvalid(m_axis_bram_58_tvalid),
        .m_axis_bram_58_tkeep(m_axis_bram_58_tkeep),
        .m_axis_bram_58_tstrb(m_axis_bram_58_tstrb),
        .m_axis_bram_58_tdata(m_axis_bram_58_tdata),
        .m_axis_bram_58_tready(m_axis_bram_58_tready),
        .ap_bram_58_addr0(ap_bram_oarg_58_addr0),
        .ap_bram_58_din0(ap_bram_oarg_58_din0),
        .ap_bram_58_dout0(ap_bram_oarg_58_dout0),
        .ap_bram_58_we0(ap_bram_oarg_58_we0),
        .ap_bram_58_en0(ap_bram_oarg_58_en0),
        .ap_bram_58_addr1(ap_bram_oarg_58_addr1),
        .ap_bram_58_din1(ap_bram_oarg_58_din1),
        .ap_bram_58_dout1(ap_bram_oarg_58_dout1),
        .ap_bram_58_we1(ap_bram_oarg_58_we1),
        .ap_bram_58_en1(ap_bram_oarg_58_en1),
        .m_axis_bram_59_tlast(m_axis_bram_59_tlast),
        .m_axis_bram_59_tvalid(m_axis_bram_59_tvalid),
        .m_axis_bram_59_tkeep(m_axis_bram_59_tkeep),
        .m_axis_bram_59_tstrb(m_axis_bram_59_tstrb),
        .m_axis_bram_59_tdata(m_axis_bram_59_tdata),
        .m_axis_bram_59_tready(m_axis_bram_59_tready),
        .ap_bram_59_addr0(ap_bram_oarg_59_addr0),
        .ap_bram_59_din0(ap_bram_oarg_59_din0),
        .ap_bram_59_dout0(ap_bram_oarg_59_dout0),
        .ap_bram_59_we0(ap_bram_oarg_59_we0),
        .ap_bram_59_en0(ap_bram_oarg_59_en0),
        .ap_bram_59_addr1(ap_bram_oarg_59_addr1),
        .ap_bram_59_din1(ap_bram_oarg_59_din1),
        .ap_bram_59_dout1(ap_bram_oarg_59_dout1),
        .ap_bram_59_we1(ap_bram_oarg_59_we1),
        .ap_bram_59_en1(ap_bram_oarg_59_en1),
        .m_axis_bram_60_tlast(m_axis_bram_60_tlast),
        .m_axis_bram_60_tvalid(m_axis_bram_60_tvalid),
        .m_axis_bram_60_tkeep(m_axis_bram_60_tkeep),
        .m_axis_bram_60_tstrb(m_axis_bram_60_tstrb),
        .m_axis_bram_60_tdata(m_axis_bram_60_tdata),
        .m_axis_bram_60_tready(m_axis_bram_60_tready),
        .ap_bram_60_addr0(ap_bram_oarg_60_addr0),
        .ap_bram_60_din0(ap_bram_oarg_60_din0),
        .ap_bram_60_dout0(ap_bram_oarg_60_dout0),
        .ap_bram_60_we0(ap_bram_oarg_60_we0),
        .ap_bram_60_en0(ap_bram_oarg_60_en0),
        .ap_bram_60_addr1(ap_bram_oarg_60_addr1),
        .ap_bram_60_din1(ap_bram_oarg_60_din1),
        .ap_bram_60_dout1(ap_bram_oarg_60_dout1),
        .ap_bram_60_we1(ap_bram_oarg_60_we1),
        .ap_bram_60_en1(ap_bram_oarg_60_en1),
        .m_axis_bram_61_tlast(m_axis_bram_61_tlast),
        .m_axis_bram_61_tvalid(m_axis_bram_61_tvalid),
        .m_axis_bram_61_tkeep(m_axis_bram_61_tkeep),
        .m_axis_bram_61_tstrb(m_axis_bram_61_tstrb),
        .m_axis_bram_61_tdata(m_axis_bram_61_tdata),
        .m_axis_bram_61_tready(m_axis_bram_61_tready),
        .ap_bram_61_addr0(ap_bram_oarg_61_addr0),
        .ap_bram_61_din0(ap_bram_oarg_61_din0),
        .ap_bram_61_dout0(ap_bram_oarg_61_dout0),
        .ap_bram_61_we0(ap_bram_oarg_61_we0),
        .ap_bram_61_en0(ap_bram_oarg_61_en0),
        .ap_bram_61_addr1(ap_bram_oarg_61_addr1),
        .ap_bram_61_din1(ap_bram_oarg_61_din1),
        .ap_bram_61_dout1(ap_bram_oarg_61_dout1),
        .ap_bram_61_we1(ap_bram_oarg_61_we1),
        .ap_bram_61_en1(ap_bram_oarg_61_en1),
        .m_axis_bram_62_tlast(m_axis_bram_62_tlast),
        .m_axis_bram_62_tvalid(m_axis_bram_62_tvalid),
        .m_axis_bram_62_tkeep(m_axis_bram_62_tkeep),
        .m_axis_bram_62_tstrb(m_axis_bram_62_tstrb),
        .m_axis_bram_62_tdata(m_axis_bram_62_tdata),
        .m_axis_bram_62_tready(m_axis_bram_62_tready),
        .ap_bram_62_addr0(ap_bram_oarg_62_addr0),
        .ap_bram_62_din0(ap_bram_oarg_62_din0),
        .ap_bram_62_dout0(ap_bram_oarg_62_dout0),
        .ap_bram_62_we0(ap_bram_oarg_62_we0),
        .ap_bram_62_en0(ap_bram_oarg_62_en0),
        .ap_bram_62_addr1(ap_bram_oarg_62_addr1),
        .ap_bram_62_din1(ap_bram_oarg_62_din1),
        .ap_bram_62_dout1(ap_bram_oarg_62_dout1),
        .ap_bram_62_we1(ap_bram_oarg_62_we1),
        .ap_bram_62_en1(ap_bram_oarg_62_en1),
        .m_axis_bram_63_tlast(m_axis_bram_63_tlast),
        .m_axis_bram_63_tvalid(m_axis_bram_63_tvalid),
        .m_axis_bram_63_tkeep(m_axis_bram_63_tkeep),
        .m_axis_bram_63_tstrb(m_axis_bram_63_tstrb),
        .m_axis_bram_63_tdata(m_axis_bram_63_tdata),
        .m_axis_bram_63_tready(m_axis_bram_63_tready),
        .ap_bram_63_addr0(ap_bram_oarg_63_addr0),
        .ap_bram_63_din0(ap_bram_oarg_63_din0),
        .ap_bram_63_dout0(ap_bram_oarg_63_dout0),
        .ap_bram_63_we0(ap_bram_oarg_63_we0),
        .ap_bram_63_en0(ap_bram_oarg_63_en0),
        .ap_bram_63_addr1(ap_bram_oarg_63_addr1),
        .ap_bram_63_din1(ap_bram_oarg_63_din1),
        .ap_bram_63_dout1(ap_bram_oarg_63_dout1),
        .ap_bram_63_we1(ap_bram_oarg_63_we1),
        .ap_bram_63_en1(ap_bram_oarg_63_en1),
        .m_axis_bram_64_tlast(m_axis_bram_64_tlast),
        .m_axis_bram_64_tvalid(m_axis_bram_64_tvalid),
        .m_axis_bram_64_tkeep(m_axis_bram_64_tkeep),
        .m_axis_bram_64_tstrb(m_axis_bram_64_tstrb),
        .m_axis_bram_64_tdata(m_axis_bram_64_tdata),
        .m_axis_bram_64_tready(m_axis_bram_64_tready),
        .ap_bram_64_addr0(ap_bram_oarg_64_addr0),
        .ap_bram_64_din0(ap_bram_oarg_64_din0),
        .ap_bram_64_dout0(ap_bram_oarg_64_dout0),
        .ap_bram_64_we0(ap_bram_oarg_64_we0),
        .ap_bram_64_en0(ap_bram_oarg_64_en0),
        .ap_bram_64_addr1(ap_bram_oarg_64_addr1),
        .ap_bram_64_din1(ap_bram_oarg_64_din1),
        .ap_bram_64_dout1(ap_bram_oarg_64_dout1),
        .ap_bram_64_we1(ap_bram_oarg_64_we1),
        .ap_bram_64_en1(ap_bram_oarg_64_en1),
        .m_axis_bram_65_tlast(m_axis_bram_65_tlast),
        .m_axis_bram_65_tvalid(m_axis_bram_65_tvalid),
        .m_axis_bram_65_tkeep(m_axis_bram_65_tkeep),
        .m_axis_bram_65_tstrb(m_axis_bram_65_tstrb),
        .m_axis_bram_65_tdata(m_axis_bram_65_tdata),
        .m_axis_bram_65_tready(m_axis_bram_65_tready),
        .ap_bram_65_addr0(ap_bram_oarg_65_addr0),
        .ap_bram_65_din0(ap_bram_oarg_65_din0),
        .ap_bram_65_dout0(ap_bram_oarg_65_dout0),
        .ap_bram_65_we0(ap_bram_oarg_65_we0),
        .ap_bram_65_en0(ap_bram_oarg_65_en0),
        .ap_bram_65_addr1(ap_bram_oarg_65_addr1),
        .ap_bram_65_din1(ap_bram_oarg_65_din1),
        .ap_bram_65_dout1(ap_bram_oarg_65_dout1),
        .ap_bram_65_we1(ap_bram_oarg_65_we1),
        .ap_bram_65_en1(ap_bram_oarg_65_en1),
        .m_axis_bram_66_tlast(m_axis_bram_66_tlast),
        .m_axis_bram_66_tvalid(m_axis_bram_66_tvalid),
        .m_axis_bram_66_tkeep(m_axis_bram_66_tkeep),
        .m_axis_bram_66_tstrb(m_axis_bram_66_tstrb),
        .m_axis_bram_66_tdata(m_axis_bram_66_tdata),
        .m_axis_bram_66_tready(m_axis_bram_66_tready),
        .ap_bram_66_addr0(ap_bram_oarg_66_addr0),
        .ap_bram_66_din0(ap_bram_oarg_66_din0),
        .ap_bram_66_dout0(ap_bram_oarg_66_dout0),
        .ap_bram_66_we0(ap_bram_oarg_66_we0),
        .ap_bram_66_en0(ap_bram_oarg_66_en0),
        .ap_bram_66_addr1(ap_bram_oarg_66_addr1),
        .ap_bram_66_din1(ap_bram_oarg_66_din1),
        .ap_bram_66_dout1(ap_bram_oarg_66_dout1),
        .ap_bram_66_we1(ap_bram_oarg_66_we1),
        .ap_bram_66_en1(ap_bram_oarg_66_en1),
        .m_axis_bram_67_tlast(m_axis_bram_67_tlast),
        .m_axis_bram_67_tvalid(m_axis_bram_67_tvalid),
        .m_axis_bram_67_tkeep(m_axis_bram_67_tkeep),
        .m_axis_bram_67_tstrb(m_axis_bram_67_tstrb),
        .m_axis_bram_67_tdata(m_axis_bram_67_tdata),
        .m_axis_bram_67_tready(m_axis_bram_67_tready),
        .ap_bram_67_addr0(ap_bram_oarg_67_addr0),
        .ap_bram_67_din0(ap_bram_oarg_67_din0),
        .ap_bram_67_dout0(ap_bram_oarg_67_dout0),
        .ap_bram_67_we0(ap_bram_oarg_67_we0),
        .ap_bram_67_en0(ap_bram_oarg_67_en0),
        .ap_bram_67_addr1(ap_bram_oarg_67_addr1),
        .ap_bram_67_din1(ap_bram_oarg_67_din1),
        .ap_bram_67_dout1(ap_bram_oarg_67_dout1),
        .ap_bram_67_we1(ap_bram_oarg_67_we1),
        .ap_bram_67_en1(ap_bram_oarg_67_en1),
        .m_axis_bram_68_tlast(m_axis_bram_68_tlast),
        .m_axis_bram_68_tvalid(m_axis_bram_68_tvalid),
        .m_axis_bram_68_tkeep(m_axis_bram_68_tkeep),
        .m_axis_bram_68_tstrb(m_axis_bram_68_tstrb),
        .m_axis_bram_68_tdata(m_axis_bram_68_tdata),
        .m_axis_bram_68_tready(m_axis_bram_68_tready),
        .ap_bram_68_addr0(ap_bram_oarg_68_addr0),
        .ap_bram_68_din0(ap_bram_oarg_68_din0),
        .ap_bram_68_dout0(ap_bram_oarg_68_dout0),
        .ap_bram_68_we0(ap_bram_oarg_68_we0),
        .ap_bram_68_en0(ap_bram_oarg_68_en0),
        .ap_bram_68_addr1(ap_bram_oarg_68_addr1),
        .ap_bram_68_din1(ap_bram_oarg_68_din1),
        .ap_bram_68_dout1(ap_bram_oarg_68_dout1),
        .ap_bram_68_we1(ap_bram_oarg_68_we1),
        .ap_bram_68_en1(ap_bram_oarg_68_en1),
        .m_axis_bram_69_tlast(m_axis_bram_69_tlast),
        .m_axis_bram_69_tvalid(m_axis_bram_69_tvalid),
        .m_axis_bram_69_tkeep(m_axis_bram_69_tkeep),
        .m_axis_bram_69_tstrb(m_axis_bram_69_tstrb),
        .m_axis_bram_69_tdata(m_axis_bram_69_tdata),
        .m_axis_bram_69_tready(m_axis_bram_69_tready),
        .ap_bram_69_addr0(ap_bram_oarg_69_addr0),
        .ap_bram_69_din0(ap_bram_oarg_69_din0),
        .ap_bram_69_dout0(ap_bram_oarg_69_dout0),
        .ap_bram_69_we0(ap_bram_oarg_69_we0),
        .ap_bram_69_en0(ap_bram_oarg_69_en0),
        .ap_bram_69_addr1(ap_bram_oarg_69_addr1),
        .ap_bram_69_din1(ap_bram_oarg_69_din1),
        .ap_bram_69_dout1(ap_bram_oarg_69_dout1),
        .ap_bram_69_we1(ap_bram_oarg_69_we1),
        .ap_bram_69_en1(ap_bram_oarg_69_en1),
        .m_axis_bram_70_tlast(m_axis_bram_70_tlast),
        .m_axis_bram_70_tvalid(m_axis_bram_70_tvalid),
        .m_axis_bram_70_tkeep(m_axis_bram_70_tkeep),
        .m_axis_bram_70_tstrb(m_axis_bram_70_tstrb),
        .m_axis_bram_70_tdata(m_axis_bram_70_tdata),
        .m_axis_bram_70_tready(m_axis_bram_70_tready),
        .ap_bram_70_addr0(ap_bram_oarg_70_addr0),
        .ap_bram_70_din0(ap_bram_oarg_70_din0),
        .ap_bram_70_dout0(ap_bram_oarg_70_dout0),
        .ap_bram_70_we0(ap_bram_oarg_70_we0),
        .ap_bram_70_en0(ap_bram_oarg_70_en0),
        .ap_bram_70_addr1(ap_bram_oarg_70_addr1),
        .ap_bram_70_din1(ap_bram_oarg_70_din1),
        .ap_bram_70_dout1(ap_bram_oarg_70_dout1),
        .ap_bram_70_we1(ap_bram_oarg_70_we1),
        .ap_bram_70_en1(ap_bram_oarg_70_en1),
        .m_axis_bram_71_tlast(m_axis_bram_71_tlast),
        .m_axis_bram_71_tvalid(m_axis_bram_71_tvalid),
        .m_axis_bram_71_tkeep(m_axis_bram_71_tkeep),
        .m_axis_bram_71_tstrb(m_axis_bram_71_tstrb),
        .m_axis_bram_71_tdata(m_axis_bram_71_tdata),
        .m_axis_bram_71_tready(m_axis_bram_71_tready),
        .ap_bram_71_addr0(ap_bram_oarg_71_addr0),
        .ap_bram_71_din0(ap_bram_oarg_71_din0),
        .ap_bram_71_dout0(ap_bram_oarg_71_dout0),
        .ap_bram_71_we0(ap_bram_oarg_71_we0),
        .ap_bram_71_en0(ap_bram_oarg_71_en0),
        .ap_bram_71_addr1(ap_bram_oarg_71_addr1),
        .ap_bram_71_din1(ap_bram_oarg_71_din1),
        .ap_bram_71_dout1(ap_bram_oarg_71_dout1),
        .ap_bram_71_we1(ap_bram_oarg_71_we1),
        .ap_bram_71_en1(ap_bram_oarg_71_en1),
        .m_axis_bram_72_tlast(m_axis_bram_72_tlast),
        .m_axis_bram_72_tvalid(m_axis_bram_72_tvalid),
        .m_axis_bram_72_tkeep(m_axis_bram_72_tkeep),
        .m_axis_bram_72_tstrb(m_axis_bram_72_tstrb),
        .m_axis_bram_72_tdata(m_axis_bram_72_tdata),
        .m_axis_bram_72_tready(m_axis_bram_72_tready),
        .ap_bram_72_addr0(ap_bram_oarg_72_addr0),
        .ap_bram_72_din0(ap_bram_oarg_72_din0),
        .ap_bram_72_dout0(ap_bram_oarg_72_dout0),
        .ap_bram_72_we0(ap_bram_oarg_72_we0),
        .ap_bram_72_en0(ap_bram_oarg_72_en0),
        .ap_bram_72_addr1(ap_bram_oarg_72_addr1),
        .ap_bram_72_din1(ap_bram_oarg_72_din1),
        .ap_bram_72_dout1(ap_bram_oarg_72_dout1),
        .ap_bram_72_we1(ap_bram_oarg_72_we1),
        .ap_bram_72_en1(ap_bram_oarg_72_en1),
        .m_axis_bram_73_tlast(m_axis_bram_73_tlast),
        .m_axis_bram_73_tvalid(m_axis_bram_73_tvalid),
        .m_axis_bram_73_tkeep(m_axis_bram_73_tkeep),
        .m_axis_bram_73_tstrb(m_axis_bram_73_tstrb),
        .m_axis_bram_73_tdata(m_axis_bram_73_tdata),
        .m_axis_bram_73_tready(m_axis_bram_73_tready),
        .ap_bram_73_addr0(ap_bram_oarg_73_addr0),
        .ap_bram_73_din0(ap_bram_oarg_73_din0),
        .ap_bram_73_dout0(ap_bram_oarg_73_dout0),
        .ap_bram_73_we0(ap_bram_oarg_73_we0),
        .ap_bram_73_en0(ap_bram_oarg_73_en0),
        .ap_bram_73_addr1(ap_bram_oarg_73_addr1),
        .ap_bram_73_din1(ap_bram_oarg_73_din1),
        .ap_bram_73_dout1(ap_bram_oarg_73_dout1),
        .ap_bram_73_we1(ap_bram_oarg_73_we1),
        .ap_bram_73_en1(ap_bram_oarg_73_en1),
        .m_axis_bram_74_tlast(m_axis_bram_74_tlast),
        .m_axis_bram_74_tvalid(m_axis_bram_74_tvalid),
        .m_axis_bram_74_tkeep(m_axis_bram_74_tkeep),
        .m_axis_bram_74_tstrb(m_axis_bram_74_tstrb),
        .m_axis_bram_74_tdata(m_axis_bram_74_tdata),
        .m_axis_bram_74_tready(m_axis_bram_74_tready),
        .ap_bram_74_addr0(ap_bram_oarg_74_addr0),
        .ap_bram_74_din0(ap_bram_oarg_74_din0),
        .ap_bram_74_dout0(ap_bram_oarg_74_dout0),
        .ap_bram_74_we0(ap_bram_oarg_74_we0),
        .ap_bram_74_en0(ap_bram_oarg_74_en0),
        .ap_bram_74_addr1(ap_bram_oarg_74_addr1),
        .ap_bram_74_din1(ap_bram_oarg_74_din1),
        .ap_bram_74_dout1(ap_bram_oarg_74_dout1),
        .ap_bram_74_we1(ap_bram_oarg_74_we1),
        .ap_bram_74_en1(ap_bram_oarg_74_en1),
        .m_axis_bram_75_tlast(m_axis_bram_75_tlast),
        .m_axis_bram_75_tvalid(m_axis_bram_75_tvalid),
        .m_axis_bram_75_tkeep(m_axis_bram_75_tkeep),
        .m_axis_bram_75_tstrb(m_axis_bram_75_tstrb),
        .m_axis_bram_75_tdata(m_axis_bram_75_tdata),
        .m_axis_bram_75_tready(m_axis_bram_75_tready),
        .ap_bram_75_addr0(ap_bram_oarg_75_addr0),
        .ap_bram_75_din0(ap_bram_oarg_75_din0),
        .ap_bram_75_dout0(ap_bram_oarg_75_dout0),
        .ap_bram_75_we0(ap_bram_oarg_75_we0),
        .ap_bram_75_en0(ap_bram_oarg_75_en0),
        .ap_bram_75_addr1(ap_bram_oarg_75_addr1),
        .ap_bram_75_din1(ap_bram_oarg_75_din1),
        .ap_bram_75_dout1(ap_bram_oarg_75_dout1),
        .ap_bram_75_we1(ap_bram_oarg_75_we1),
        .ap_bram_75_en1(ap_bram_oarg_75_en1),
        .m_axis_bram_76_tlast(m_axis_bram_76_tlast),
        .m_axis_bram_76_tvalid(m_axis_bram_76_tvalid),
        .m_axis_bram_76_tkeep(m_axis_bram_76_tkeep),
        .m_axis_bram_76_tstrb(m_axis_bram_76_tstrb),
        .m_axis_bram_76_tdata(m_axis_bram_76_tdata),
        .m_axis_bram_76_tready(m_axis_bram_76_tready),
        .ap_bram_76_addr0(ap_bram_oarg_76_addr0),
        .ap_bram_76_din0(ap_bram_oarg_76_din0),
        .ap_bram_76_dout0(ap_bram_oarg_76_dout0),
        .ap_bram_76_we0(ap_bram_oarg_76_we0),
        .ap_bram_76_en0(ap_bram_oarg_76_en0),
        .ap_bram_76_addr1(ap_bram_oarg_76_addr1),
        .ap_bram_76_din1(ap_bram_oarg_76_din1),
        .ap_bram_76_dout1(ap_bram_oarg_76_dout1),
        .ap_bram_76_we1(ap_bram_oarg_76_we1),
        .ap_bram_76_en1(ap_bram_oarg_76_en1),
        .m_axis_bram_77_tlast(m_axis_bram_77_tlast),
        .m_axis_bram_77_tvalid(m_axis_bram_77_tvalid),
        .m_axis_bram_77_tkeep(m_axis_bram_77_tkeep),
        .m_axis_bram_77_tstrb(m_axis_bram_77_tstrb),
        .m_axis_bram_77_tdata(m_axis_bram_77_tdata),
        .m_axis_bram_77_tready(m_axis_bram_77_tready),
        .ap_bram_77_addr0(ap_bram_oarg_77_addr0),
        .ap_bram_77_din0(ap_bram_oarg_77_din0),
        .ap_bram_77_dout0(ap_bram_oarg_77_dout0),
        .ap_bram_77_we0(ap_bram_oarg_77_we0),
        .ap_bram_77_en0(ap_bram_oarg_77_en0),
        .ap_bram_77_addr1(ap_bram_oarg_77_addr1),
        .ap_bram_77_din1(ap_bram_oarg_77_din1),
        .ap_bram_77_dout1(ap_bram_oarg_77_dout1),
        .ap_bram_77_we1(ap_bram_oarg_77_we1),
        .ap_bram_77_en1(ap_bram_oarg_77_en1),
        .m_axis_bram_78_tlast(m_axis_bram_78_tlast),
        .m_axis_bram_78_tvalid(m_axis_bram_78_tvalid),
        .m_axis_bram_78_tkeep(m_axis_bram_78_tkeep),
        .m_axis_bram_78_tstrb(m_axis_bram_78_tstrb),
        .m_axis_bram_78_tdata(m_axis_bram_78_tdata),
        .m_axis_bram_78_tready(m_axis_bram_78_tready),
        .ap_bram_78_addr0(ap_bram_oarg_78_addr0),
        .ap_bram_78_din0(ap_bram_oarg_78_din0),
        .ap_bram_78_dout0(ap_bram_oarg_78_dout0),
        .ap_bram_78_we0(ap_bram_oarg_78_we0),
        .ap_bram_78_en0(ap_bram_oarg_78_en0),
        .ap_bram_78_addr1(ap_bram_oarg_78_addr1),
        .ap_bram_78_din1(ap_bram_oarg_78_din1),
        .ap_bram_78_dout1(ap_bram_oarg_78_dout1),
        .ap_bram_78_we1(ap_bram_oarg_78_we1),
        .ap_bram_78_en1(ap_bram_oarg_78_en1),
        .m_axis_bram_79_tlast(m_axis_bram_79_tlast),
        .m_axis_bram_79_tvalid(m_axis_bram_79_tvalid),
        .m_axis_bram_79_tkeep(m_axis_bram_79_tkeep),
        .m_axis_bram_79_tstrb(m_axis_bram_79_tstrb),
        .m_axis_bram_79_tdata(m_axis_bram_79_tdata),
        .m_axis_bram_79_tready(m_axis_bram_79_tready),
        .ap_bram_79_addr0(ap_bram_oarg_79_addr0),
        .ap_bram_79_din0(ap_bram_oarg_79_din0),
        .ap_bram_79_dout0(ap_bram_oarg_79_dout0),
        .ap_bram_79_we0(ap_bram_oarg_79_we0),
        .ap_bram_79_en0(ap_bram_oarg_79_en0),
        .ap_bram_79_addr1(ap_bram_oarg_79_addr1),
        .ap_bram_79_din1(ap_bram_oarg_79_din1),
        .ap_bram_79_dout1(ap_bram_oarg_79_dout1),
        .ap_bram_79_we1(ap_bram_oarg_79_we1),
        .ap_bram_79_en1(ap_bram_oarg_79_en1),
        .m_axis_bram_80_tlast(m_axis_bram_80_tlast),
        .m_axis_bram_80_tvalid(m_axis_bram_80_tvalid),
        .m_axis_bram_80_tkeep(m_axis_bram_80_tkeep),
        .m_axis_bram_80_tstrb(m_axis_bram_80_tstrb),
        .m_axis_bram_80_tdata(m_axis_bram_80_tdata),
        .m_axis_bram_80_tready(m_axis_bram_80_tready),
        .ap_bram_80_addr0(ap_bram_oarg_80_addr0),
        .ap_bram_80_din0(ap_bram_oarg_80_din0),
        .ap_bram_80_dout0(ap_bram_oarg_80_dout0),
        .ap_bram_80_we0(ap_bram_oarg_80_we0),
        .ap_bram_80_en0(ap_bram_oarg_80_en0),
        .ap_bram_80_addr1(ap_bram_oarg_80_addr1),
        .ap_bram_80_din1(ap_bram_oarg_80_din1),
        .ap_bram_80_dout1(ap_bram_oarg_80_dout1),
        .ap_bram_80_we1(ap_bram_oarg_80_we1),
        .ap_bram_80_en1(ap_bram_oarg_80_en1),
        .m_axis_bram_81_tlast(m_axis_bram_81_tlast),
        .m_axis_bram_81_tvalid(m_axis_bram_81_tvalid),
        .m_axis_bram_81_tkeep(m_axis_bram_81_tkeep),
        .m_axis_bram_81_tstrb(m_axis_bram_81_tstrb),
        .m_axis_bram_81_tdata(m_axis_bram_81_tdata),
        .m_axis_bram_81_tready(m_axis_bram_81_tready),
        .ap_bram_81_addr0(ap_bram_oarg_81_addr0),
        .ap_bram_81_din0(ap_bram_oarg_81_din0),
        .ap_bram_81_dout0(ap_bram_oarg_81_dout0),
        .ap_bram_81_we0(ap_bram_oarg_81_we0),
        .ap_bram_81_en0(ap_bram_oarg_81_en0),
        .ap_bram_81_addr1(ap_bram_oarg_81_addr1),
        .ap_bram_81_din1(ap_bram_oarg_81_din1),
        .ap_bram_81_dout1(ap_bram_oarg_81_dout1),
        .ap_bram_81_we1(ap_bram_oarg_81_we1),
        .ap_bram_81_en1(ap_bram_oarg_81_en1),
        .m_axis_bram_82_tlast(m_axis_bram_82_tlast),
        .m_axis_bram_82_tvalid(m_axis_bram_82_tvalid),
        .m_axis_bram_82_tkeep(m_axis_bram_82_tkeep),
        .m_axis_bram_82_tstrb(m_axis_bram_82_tstrb),
        .m_axis_bram_82_tdata(m_axis_bram_82_tdata),
        .m_axis_bram_82_tready(m_axis_bram_82_tready),
        .ap_bram_82_addr0(ap_bram_oarg_82_addr0),
        .ap_bram_82_din0(ap_bram_oarg_82_din0),
        .ap_bram_82_dout0(ap_bram_oarg_82_dout0),
        .ap_bram_82_we0(ap_bram_oarg_82_we0),
        .ap_bram_82_en0(ap_bram_oarg_82_en0),
        .ap_bram_82_addr1(ap_bram_oarg_82_addr1),
        .ap_bram_82_din1(ap_bram_oarg_82_din1),
        .ap_bram_82_dout1(ap_bram_oarg_82_dout1),
        .ap_bram_82_we1(ap_bram_oarg_82_we1),
        .ap_bram_82_en1(ap_bram_oarg_82_en1),
        .m_axis_bram_83_tlast(m_axis_bram_83_tlast),
        .m_axis_bram_83_tvalid(m_axis_bram_83_tvalid),
        .m_axis_bram_83_tkeep(m_axis_bram_83_tkeep),
        .m_axis_bram_83_tstrb(m_axis_bram_83_tstrb),
        .m_axis_bram_83_tdata(m_axis_bram_83_tdata),
        .m_axis_bram_83_tready(m_axis_bram_83_tready),
        .ap_bram_83_addr0(ap_bram_oarg_83_addr0),
        .ap_bram_83_din0(ap_bram_oarg_83_din0),
        .ap_bram_83_dout0(ap_bram_oarg_83_dout0),
        .ap_bram_83_we0(ap_bram_oarg_83_we0),
        .ap_bram_83_en0(ap_bram_oarg_83_en0),
        .ap_bram_83_addr1(ap_bram_oarg_83_addr1),
        .ap_bram_83_din1(ap_bram_oarg_83_din1),
        .ap_bram_83_dout1(ap_bram_oarg_83_dout1),
        .ap_bram_83_we1(ap_bram_oarg_83_we1),
        .ap_bram_83_en1(ap_bram_oarg_83_en1),
        .m_axis_bram_84_tlast(m_axis_bram_84_tlast),
        .m_axis_bram_84_tvalid(m_axis_bram_84_tvalid),
        .m_axis_bram_84_tkeep(m_axis_bram_84_tkeep),
        .m_axis_bram_84_tstrb(m_axis_bram_84_tstrb),
        .m_axis_bram_84_tdata(m_axis_bram_84_tdata),
        .m_axis_bram_84_tready(m_axis_bram_84_tready),
        .ap_bram_84_addr0(ap_bram_oarg_84_addr0),
        .ap_bram_84_din0(ap_bram_oarg_84_din0),
        .ap_bram_84_dout0(ap_bram_oarg_84_dout0),
        .ap_bram_84_we0(ap_bram_oarg_84_we0),
        .ap_bram_84_en0(ap_bram_oarg_84_en0),
        .ap_bram_84_addr1(ap_bram_oarg_84_addr1),
        .ap_bram_84_din1(ap_bram_oarg_84_din1),
        .ap_bram_84_dout1(ap_bram_oarg_84_dout1),
        .ap_bram_84_we1(ap_bram_oarg_84_we1),
        .ap_bram_84_en1(ap_bram_oarg_84_en1),
        .m_axis_bram_85_tlast(m_axis_bram_85_tlast),
        .m_axis_bram_85_tvalid(m_axis_bram_85_tvalid),
        .m_axis_bram_85_tkeep(m_axis_bram_85_tkeep),
        .m_axis_bram_85_tstrb(m_axis_bram_85_tstrb),
        .m_axis_bram_85_tdata(m_axis_bram_85_tdata),
        .m_axis_bram_85_tready(m_axis_bram_85_tready),
        .ap_bram_85_addr0(ap_bram_oarg_85_addr0),
        .ap_bram_85_din0(ap_bram_oarg_85_din0),
        .ap_bram_85_dout0(ap_bram_oarg_85_dout0),
        .ap_bram_85_we0(ap_bram_oarg_85_we0),
        .ap_bram_85_en0(ap_bram_oarg_85_en0),
        .ap_bram_85_addr1(ap_bram_oarg_85_addr1),
        .ap_bram_85_din1(ap_bram_oarg_85_din1),
        .ap_bram_85_dout1(ap_bram_oarg_85_dout1),
        .ap_bram_85_we1(ap_bram_oarg_85_we1),
        .ap_bram_85_en1(ap_bram_oarg_85_en1),
        .m_axis_bram_86_tlast(m_axis_bram_86_tlast),
        .m_axis_bram_86_tvalid(m_axis_bram_86_tvalid),
        .m_axis_bram_86_tkeep(m_axis_bram_86_tkeep),
        .m_axis_bram_86_tstrb(m_axis_bram_86_tstrb),
        .m_axis_bram_86_tdata(m_axis_bram_86_tdata),
        .m_axis_bram_86_tready(m_axis_bram_86_tready),
        .ap_bram_86_addr0(ap_bram_oarg_86_addr0),
        .ap_bram_86_din0(ap_bram_oarg_86_din0),
        .ap_bram_86_dout0(ap_bram_oarg_86_dout0),
        .ap_bram_86_we0(ap_bram_oarg_86_we0),
        .ap_bram_86_en0(ap_bram_oarg_86_en0),
        .ap_bram_86_addr1(ap_bram_oarg_86_addr1),
        .ap_bram_86_din1(ap_bram_oarg_86_din1),
        .ap_bram_86_dout1(ap_bram_oarg_86_dout1),
        .ap_bram_86_we1(ap_bram_oarg_86_we1),
        .ap_bram_86_en1(ap_bram_oarg_86_en1),
        .m_axis_bram_87_tlast(m_axis_bram_87_tlast),
        .m_axis_bram_87_tvalid(m_axis_bram_87_tvalid),
        .m_axis_bram_87_tkeep(m_axis_bram_87_tkeep),
        .m_axis_bram_87_tstrb(m_axis_bram_87_tstrb),
        .m_axis_bram_87_tdata(m_axis_bram_87_tdata),
        .m_axis_bram_87_tready(m_axis_bram_87_tready),
        .ap_bram_87_addr0(ap_bram_oarg_87_addr0),
        .ap_bram_87_din0(ap_bram_oarg_87_din0),
        .ap_bram_87_dout0(ap_bram_oarg_87_dout0),
        .ap_bram_87_we0(ap_bram_oarg_87_we0),
        .ap_bram_87_en0(ap_bram_oarg_87_en0),
        .ap_bram_87_addr1(ap_bram_oarg_87_addr1),
        .ap_bram_87_din1(ap_bram_oarg_87_din1),
        .ap_bram_87_dout1(ap_bram_oarg_87_dout1),
        .ap_bram_87_we1(ap_bram_oarg_87_we1),
        .ap_bram_87_en1(ap_bram_oarg_87_en1),
        .m_axis_bram_88_tlast(m_axis_bram_88_tlast),
        .m_axis_bram_88_tvalid(m_axis_bram_88_tvalid),
        .m_axis_bram_88_tkeep(m_axis_bram_88_tkeep),
        .m_axis_bram_88_tstrb(m_axis_bram_88_tstrb),
        .m_axis_bram_88_tdata(m_axis_bram_88_tdata),
        .m_axis_bram_88_tready(m_axis_bram_88_tready),
        .ap_bram_88_addr0(ap_bram_oarg_88_addr0),
        .ap_bram_88_din0(ap_bram_oarg_88_din0),
        .ap_bram_88_dout0(ap_bram_oarg_88_dout0),
        .ap_bram_88_we0(ap_bram_oarg_88_we0),
        .ap_bram_88_en0(ap_bram_oarg_88_en0),
        .ap_bram_88_addr1(ap_bram_oarg_88_addr1),
        .ap_bram_88_din1(ap_bram_oarg_88_din1),
        .ap_bram_88_dout1(ap_bram_oarg_88_dout1),
        .ap_bram_88_we1(ap_bram_oarg_88_we1),
        .ap_bram_88_en1(ap_bram_oarg_88_en1),
        .m_axis_bram_89_tlast(m_axis_bram_89_tlast),
        .m_axis_bram_89_tvalid(m_axis_bram_89_tvalid),
        .m_axis_bram_89_tkeep(m_axis_bram_89_tkeep),
        .m_axis_bram_89_tstrb(m_axis_bram_89_tstrb),
        .m_axis_bram_89_tdata(m_axis_bram_89_tdata),
        .m_axis_bram_89_tready(m_axis_bram_89_tready),
        .ap_bram_89_addr0(ap_bram_oarg_89_addr0),
        .ap_bram_89_din0(ap_bram_oarg_89_din0),
        .ap_bram_89_dout0(ap_bram_oarg_89_dout0),
        .ap_bram_89_we0(ap_bram_oarg_89_we0),
        .ap_bram_89_en0(ap_bram_oarg_89_en0),
        .ap_bram_89_addr1(ap_bram_oarg_89_addr1),
        .ap_bram_89_din1(ap_bram_oarg_89_din1),
        .ap_bram_89_dout1(ap_bram_oarg_89_dout1),
        .ap_bram_89_we1(ap_bram_oarg_89_we1),
        .ap_bram_89_en1(ap_bram_oarg_89_en1),
        .m_axis_bram_90_tlast(m_axis_bram_90_tlast),
        .m_axis_bram_90_tvalid(m_axis_bram_90_tvalid),
        .m_axis_bram_90_tkeep(m_axis_bram_90_tkeep),
        .m_axis_bram_90_tstrb(m_axis_bram_90_tstrb),
        .m_axis_bram_90_tdata(m_axis_bram_90_tdata),
        .m_axis_bram_90_tready(m_axis_bram_90_tready),
        .ap_bram_90_addr0(ap_bram_oarg_90_addr0),
        .ap_bram_90_din0(ap_bram_oarg_90_din0),
        .ap_bram_90_dout0(ap_bram_oarg_90_dout0),
        .ap_bram_90_we0(ap_bram_oarg_90_we0),
        .ap_bram_90_en0(ap_bram_oarg_90_en0),
        .ap_bram_90_addr1(ap_bram_oarg_90_addr1),
        .ap_bram_90_din1(ap_bram_oarg_90_din1),
        .ap_bram_90_dout1(ap_bram_oarg_90_dout1),
        .ap_bram_90_we1(ap_bram_oarg_90_we1),
        .ap_bram_90_en1(ap_bram_oarg_90_en1),
        .m_axis_bram_91_tlast(m_axis_bram_91_tlast),
        .m_axis_bram_91_tvalid(m_axis_bram_91_tvalid),
        .m_axis_bram_91_tkeep(m_axis_bram_91_tkeep),
        .m_axis_bram_91_tstrb(m_axis_bram_91_tstrb),
        .m_axis_bram_91_tdata(m_axis_bram_91_tdata),
        .m_axis_bram_91_tready(m_axis_bram_91_tready),
        .ap_bram_91_addr0(ap_bram_oarg_91_addr0),
        .ap_bram_91_din0(ap_bram_oarg_91_din0),
        .ap_bram_91_dout0(ap_bram_oarg_91_dout0),
        .ap_bram_91_we0(ap_bram_oarg_91_we0),
        .ap_bram_91_en0(ap_bram_oarg_91_en0),
        .ap_bram_91_addr1(ap_bram_oarg_91_addr1),
        .ap_bram_91_din1(ap_bram_oarg_91_din1),
        .ap_bram_91_dout1(ap_bram_oarg_91_dout1),
        .ap_bram_91_we1(ap_bram_oarg_91_we1),
        .ap_bram_91_en1(ap_bram_oarg_91_en1),
        .m_axis_bram_92_tlast(m_axis_bram_92_tlast),
        .m_axis_bram_92_tvalid(m_axis_bram_92_tvalid),
        .m_axis_bram_92_tkeep(m_axis_bram_92_tkeep),
        .m_axis_bram_92_tstrb(m_axis_bram_92_tstrb),
        .m_axis_bram_92_tdata(m_axis_bram_92_tdata),
        .m_axis_bram_92_tready(m_axis_bram_92_tready),
        .ap_bram_92_addr0(ap_bram_oarg_92_addr0),
        .ap_bram_92_din0(ap_bram_oarg_92_din0),
        .ap_bram_92_dout0(ap_bram_oarg_92_dout0),
        .ap_bram_92_we0(ap_bram_oarg_92_we0),
        .ap_bram_92_en0(ap_bram_oarg_92_en0),
        .ap_bram_92_addr1(ap_bram_oarg_92_addr1),
        .ap_bram_92_din1(ap_bram_oarg_92_din1),
        .ap_bram_92_dout1(ap_bram_oarg_92_dout1),
        .ap_bram_92_we1(ap_bram_oarg_92_we1),
        .ap_bram_92_en1(ap_bram_oarg_92_en1),
        .m_axis_bram_93_tlast(m_axis_bram_93_tlast),
        .m_axis_bram_93_tvalid(m_axis_bram_93_tvalid),
        .m_axis_bram_93_tkeep(m_axis_bram_93_tkeep),
        .m_axis_bram_93_tstrb(m_axis_bram_93_tstrb),
        .m_axis_bram_93_tdata(m_axis_bram_93_tdata),
        .m_axis_bram_93_tready(m_axis_bram_93_tready),
        .ap_bram_93_addr0(ap_bram_oarg_93_addr0),
        .ap_bram_93_din0(ap_bram_oarg_93_din0),
        .ap_bram_93_dout0(ap_bram_oarg_93_dout0),
        .ap_bram_93_we0(ap_bram_oarg_93_we0),
        .ap_bram_93_en0(ap_bram_oarg_93_en0),
        .ap_bram_93_addr1(ap_bram_oarg_93_addr1),
        .ap_bram_93_din1(ap_bram_oarg_93_din1),
        .ap_bram_93_dout1(ap_bram_oarg_93_dout1),
        .ap_bram_93_we1(ap_bram_oarg_93_we1),
        .ap_bram_93_en1(ap_bram_oarg_93_en1),
        .m_axis_bram_94_tlast(m_axis_bram_94_tlast),
        .m_axis_bram_94_tvalid(m_axis_bram_94_tvalid),
        .m_axis_bram_94_tkeep(m_axis_bram_94_tkeep),
        .m_axis_bram_94_tstrb(m_axis_bram_94_tstrb),
        .m_axis_bram_94_tdata(m_axis_bram_94_tdata),
        .m_axis_bram_94_tready(m_axis_bram_94_tready),
        .ap_bram_94_addr0(ap_bram_oarg_94_addr0),
        .ap_bram_94_din0(ap_bram_oarg_94_din0),
        .ap_bram_94_dout0(ap_bram_oarg_94_dout0),
        .ap_bram_94_we0(ap_bram_oarg_94_we0),
        .ap_bram_94_en0(ap_bram_oarg_94_en0),
        .ap_bram_94_addr1(ap_bram_oarg_94_addr1),
        .ap_bram_94_din1(ap_bram_oarg_94_din1),
        .ap_bram_94_dout1(ap_bram_oarg_94_dout1),
        .ap_bram_94_we1(ap_bram_oarg_94_we1),
        .ap_bram_94_en1(ap_bram_oarg_94_en1),
        .m_axis_bram_95_tlast(m_axis_bram_95_tlast),
        .m_axis_bram_95_tvalid(m_axis_bram_95_tvalid),
        .m_axis_bram_95_tkeep(m_axis_bram_95_tkeep),
        .m_axis_bram_95_tstrb(m_axis_bram_95_tstrb),
        .m_axis_bram_95_tdata(m_axis_bram_95_tdata),
        .m_axis_bram_95_tready(m_axis_bram_95_tready),
        .ap_bram_95_addr0(ap_bram_oarg_95_addr0),
        .ap_bram_95_din0(ap_bram_oarg_95_din0),
        .ap_bram_95_dout0(ap_bram_oarg_95_dout0),
        .ap_bram_95_we0(ap_bram_oarg_95_we0),
        .ap_bram_95_en0(ap_bram_oarg_95_en0),
        .ap_bram_95_addr1(ap_bram_oarg_95_addr1),
        .ap_bram_95_din1(ap_bram_oarg_95_din1),
        .ap_bram_95_dout1(ap_bram_oarg_95_dout1),
        .ap_bram_95_we1(ap_bram_oarg_95_we1),
        .ap_bram_95_en1(ap_bram_oarg_95_en1),
        .m_axis_bram_96_tlast(m_axis_bram_96_tlast),
        .m_axis_bram_96_tvalid(m_axis_bram_96_tvalid),
        .m_axis_bram_96_tkeep(m_axis_bram_96_tkeep),
        .m_axis_bram_96_tstrb(m_axis_bram_96_tstrb),
        .m_axis_bram_96_tdata(m_axis_bram_96_tdata),
        .m_axis_bram_96_tready(m_axis_bram_96_tready),
        .ap_bram_96_addr0(ap_bram_oarg_96_addr0),
        .ap_bram_96_din0(ap_bram_oarg_96_din0),
        .ap_bram_96_dout0(ap_bram_oarg_96_dout0),
        .ap_bram_96_we0(ap_bram_oarg_96_we0),
        .ap_bram_96_en0(ap_bram_oarg_96_en0),
        .ap_bram_96_addr1(ap_bram_oarg_96_addr1),
        .ap_bram_96_din1(ap_bram_oarg_96_din1),
        .ap_bram_96_dout1(ap_bram_oarg_96_dout1),
        .ap_bram_96_we1(ap_bram_oarg_96_we1),
        .ap_bram_96_en1(ap_bram_oarg_96_en1),
        .m_axis_bram_97_tlast(m_axis_bram_97_tlast),
        .m_axis_bram_97_tvalid(m_axis_bram_97_tvalid),
        .m_axis_bram_97_tkeep(m_axis_bram_97_tkeep),
        .m_axis_bram_97_tstrb(m_axis_bram_97_tstrb),
        .m_axis_bram_97_tdata(m_axis_bram_97_tdata),
        .m_axis_bram_97_tready(m_axis_bram_97_tready),
        .ap_bram_97_addr0(ap_bram_oarg_97_addr0),
        .ap_bram_97_din0(ap_bram_oarg_97_din0),
        .ap_bram_97_dout0(ap_bram_oarg_97_dout0),
        .ap_bram_97_we0(ap_bram_oarg_97_we0),
        .ap_bram_97_en0(ap_bram_oarg_97_en0),
        .ap_bram_97_addr1(ap_bram_oarg_97_addr1),
        .ap_bram_97_din1(ap_bram_oarg_97_din1),
        .ap_bram_97_dout1(ap_bram_oarg_97_dout1),
        .ap_bram_97_we1(ap_bram_oarg_97_we1),
        .ap_bram_97_en1(ap_bram_oarg_97_en1),
        .m_axis_bram_98_tlast(m_axis_bram_98_tlast),
        .m_axis_bram_98_tvalid(m_axis_bram_98_tvalid),
        .m_axis_bram_98_tkeep(m_axis_bram_98_tkeep),
        .m_axis_bram_98_tstrb(m_axis_bram_98_tstrb),
        .m_axis_bram_98_tdata(m_axis_bram_98_tdata),
        .m_axis_bram_98_tready(m_axis_bram_98_tready),
        .ap_bram_98_addr0(ap_bram_oarg_98_addr0),
        .ap_bram_98_din0(ap_bram_oarg_98_din0),
        .ap_bram_98_dout0(ap_bram_oarg_98_dout0),
        .ap_bram_98_we0(ap_bram_oarg_98_we0),
        .ap_bram_98_en0(ap_bram_oarg_98_en0),
        .ap_bram_98_addr1(ap_bram_oarg_98_addr1),
        .ap_bram_98_din1(ap_bram_oarg_98_din1),
        .ap_bram_98_dout1(ap_bram_oarg_98_dout1),
        .ap_bram_98_we1(ap_bram_oarg_98_we1),
        .ap_bram_98_en1(ap_bram_oarg_98_en1),
        .m_axis_bram_99_tlast(m_axis_bram_99_tlast),
        .m_axis_bram_99_tvalid(m_axis_bram_99_tvalid),
        .m_axis_bram_99_tkeep(m_axis_bram_99_tkeep),
        .m_axis_bram_99_tstrb(m_axis_bram_99_tstrb),
        .m_axis_bram_99_tdata(m_axis_bram_99_tdata),
        .m_axis_bram_99_tready(m_axis_bram_99_tready),
        .ap_bram_99_addr0(ap_bram_oarg_99_addr0),
        .ap_bram_99_din0(ap_bram_oarg_99_din0),
        .ap_bram_99_dout0(ap_bram_oarg_99_dout0),
        .ap_bram_99_we0(ap_bram_oarg_99_we0),
        .ap_bram_99_en0(ap_bram_oarg_99_en0),
        .ap_bram_99_addr1(ap_bram_oarg_99_addr1),
        .ap_bram_99_din1(ap_bram_oarg_99_din1),
        .ap_bram_99_dout1(ap_bram_oarg_99_dout1),
        .ap_bram_99_we1(ap_bram_oarg_99_we1),
        .ap_bram_99_en1(ap_bram_oarg_99_en1),
        .m_axis_bram_100_tlast(m_axis_bram_100_tlast),
        .m_axis_bram_100_tvalid(m_axis_bram_100_tvalid),
        .m_axis_bram_100_tkeep(m_axis_bram_100_tkeep),
        .m_axis_bram_100_tstrb(m_axis_bram_100_tstrb),
        .m_axis_bram_100_tdata(m_axis_bram_100_tdata),
        .m_axis_bram_100_tready(m_axis_bram_100_tready),
        .ap_bram_100_addr0(ap_bram_oarg_100_addr0),
        .ap_bram_100_din0(ap_bram_oarg_100_din0),
        .ap_bram_100_dout0(ap_bram_oarg_100_dout0),
        .ap_bram_100_we0(ap_bram_oarg_100_we0),
        .ap_bram_100_en0(ap_bram_oarg_100_en0),
        .ap_bram_100_addr1(ap_bram_oarg_100_addr1),
        .ap_bram_100_din1(ap_bram_oarg_100_din1),
        .ap_bram_100_dout1(ap_bram_oarg_100_dout1),
        .ap_bram_100_we1(ap_bram_oarg_100_we1),
        .ap_bram_100_en1(ap_bram_oarg_100_en1),
        .m_axis_bram_101_tlast(m_axis_bram_101_tlast),
        .m_axis_bram_101_tvalid(m_axis_bram_101_tvalid),
        .m_axis_bram_101_tkeep(m_axis_bram_101_tkeep),
        .m_axis_bram_101_tstrb(m_axis_bram_101_tstrb),
        .m_axis_bram_101_tdata(m_axis_bram_101_tdata),
        .m_axis_bram_101_tready(m_axis_bram_101_tready),
        .ap_bram_101_addr0(ap_bram_oarg_101_addr0),
        .ap_bram_101_din0(ap_bram_oarg_101_din0),
        .ap_bram_101_dout0(ap_bram_oarg_101_dout0),
        .ap_bram_101_we0(ap_bram_oarg_101_we0),
        .ap_bram_101_en0(ap_bram_oarg_101_en0),
        .ap_bram_101_addr1(ap_bram_oarg_101_addr1),
        .ap_bram_101_din1(ap_bram_oarg_101_din1),
        .ap_bram_101_dout1(ap_bram_oarg_101_dout1),
        .ap_bram_101_we1(ap_bram_oarg_101_we1),
        .ap_bram_101_en1(ap_bram_oarg_101_en1),
        .m_axis_bram_102_tlast(m_axis_bram_102_tlast),
        .m_axis_bram_102_tvalid(m_axis_bram_102_tvalid),
        .m_axis_bram_102_tkeep(m_axis_bram_102_tkeep),
        .m_axis_bram_102_tstrb(m_axis_bram_102_tstrb),
        .m_axis_bram_102_tdata(m_axis_bram_102_tdata),
        .m_axis_bram_102_tready(m_axis_bram_102_tready),
        .ap_bram_102_addr0(ap_bram_oarg_102_addr0),
        .ap_bram_102_din0(ap_bram_oarg_102_din0),
        .ap_bram_102_dout0(ap_bram_oarg_102_dout0),
        .ap_bram_102_we0(ap_bram_oarg_102_we0),
        .ap_bram_102_en0(ap_bram_oarg_102_en0),
        .ap_bram_102_addr1(ap_bram_oarg_102_addr1),
        .ap_bram_102_din1(ap_bram_oarg_102_din1),
        .ap_bram_102_dout1(ap_bram_oarg_102_dout1),
        .ap_bram_102_we1(ap_bram_oarg_102_we1),
        .ap_bram_102_en1(ap_bram_oarg_102_en1),
        .m_axis_bram_103_tlast(m_axis_bram_103_tlast),
        .m_axis_bram_103_tvalid(m_axis_bram_103_tvalid),
        .m_axis_bram_103_tkeep(m_axis_bram_103_tkeep),
        .m_axis_bram_103_tstrb(m_axis_bram_103_tstrb),
        .m_axis_bram_103_tdata(m_axis_bram_103_tdata),
        .m_axis_bram_103_tready(m_axis_bram_103_tready),
        .ap_bram_103_addr0(ap_bram_oarg_103_addr0),
        .ap_bram_103_din0(ap_bram_oarg_103_din0),
        .ap_bram_103_dout0(ap_bram_oarg_103_dout0),
        .ap_bram_103_we0(ap_bram_oarg_103_we0),
        .ap_bram_103_en0(ap_bram_oarg_103_en0),
        .ap_bram_103_addr1(ap_bram_oarg_103_addr1),
        .ap_bram_103_din1(ap_bram_oarg_103_din1),
        .ap_bram_103_dout1(ap_bram_oarg_103_dout1),
        .ap_bram_103_we1(ap_bram_oarg_103_we1),
        .ap_bram_103_en1(ap_bram_oarg_103_en1),
        .m_axis_bram_104_tlast(m_axis_bram_104_tlast),
        .m_axis_bram_104_tvalid(m_axis_bram_104_tvalid),
        .m_axis_bram_104_tkeep(m_axis_bram_104_tkeep),
        .m_axis_bram_104_tstrb(m_axis_bram_104_tstrb),
        .m_axis_bram_104_tdata(m_axis_bram_104_tdata),
        .m_axis_bram_104_tready(m_axis_bram_104_tready),
        .ap_bram_104_addr0(ap_bram_oarg_104_addr0),
        .ap_bram_104_din0(ap_bram_oarg_104_din0),
        .ap_bram_104_dout0(ap_bram_oarg_104_dout0),
        .ap_bram_104_we0(ap_bram_oarg_104_we0),
        .ap_bram_104_en0(ap_bram_oarg_104_en0),
        .ap_bram_104_addr1(ap_bram_oarg_104_addr1),
        .ap_bram_104_din1(ap_bram_oarg_104_din1),
        .ap_bram_104_dout1(ap_bram_oarg_104_dout1),
        .ap_bram_104_we1(ap_bram_oarg_104_we1),
        .ap_bram_104_en1(ap_bram_oarg_104_en1),
        .m_axis_bram_105_tlast(m_axis_bram_105_tlast),
        .m_axis_bram_105_tvalid(m_axis_bram_105_tvalid),
        .m_axis_bram_105_tkeep(m_axis_bram_105_tkeep),
        .m_axis_bram_105_tstrb(m_axis_bram_105_tstrb),
        .m_axis_bram_105_tdata(m_axis_bram_105_tdata),
        .m_axis_bram_105_tready(m_axis_bram_105_tready),
        .ap_bram_105_addr0(ap_bram_oarg_105_addr0),
        .ap_bram_105_din0(ap_bram_oarg_105_din0),
        .ap_bram_105_dout0(ap_bram_oarg_105_dout0),
        .ap_bram_105_we0(ap_bram_oarg_105_we0),
        .ap_bram_105_en0(ap_bram_oarg_105_en0),
        .ap_bram_105_addr1(ap_bram_oarg_105_addr1),
        .ap_bram_105_din1(ap_bram_oarg_105_din1),
        .ap_bram_105_dout1(ap_bram_oarg_105_dout1),
        .ap_bram_105_we1(ap_bram_oarg_105_we1),
        .ap_bram_105_en1(ap_bram_oarg_105_en1),
        .m_axis_bram_106_tlast(m_axis_bram_106_tlast),
        .m_axis_bram_106_tvalid(m_axis_bram_106_tvalid),
        .m_axis_bram_106_tkeep(m_axis_bram_106_tkeep),
        .m_axis_bram_106_tstrb(m_axis_bram_106_tstrb),
        .m_axis_bram_106_tdata(m_axis_bram_106_tdata),
        .m_axis_bram_106_tready(m_axis_bram_106_tready),
        .ap_bram_106_addr0(ap_bram_oarg_106_addr0),
        .ap_bram_106_din0(ap_bram_oarg_106_din0),
        .ap_bram_106_dout0(ap_bram_oarg_106_dout0),
        .ap_bram_106_we0(ap_bram_oarg_106_we0),
        .ap_bram_106_en0(ap_bram_oarg_106_en0),
        .ap_bram_106_addr1(ap_bram_oarg_106_addr1),
        .ap_bram_106_din1(ap_bram_oarg_106_din1),
        .ap_bram_106_dout1(ap_bram_oarg_106_dout1),
        .ap_bram_106_we1(ap_bram_oarg_106_we1),
        .ap_bram_106_en1(ap_bram_oarg_106_en1),
        .m_axis_bram_107_tlast(m_axis_bram_107_tlast),
        .m_axis_bram_107_tvalid(m_axis_bram_107_tvalid),
        .m_axis_bram_107_tkeep(m_axis_bram_107_tkeep),
        .m_axis_bram_107_tstrb(m_axis_bram_107_tstrb),
        .m_axis_bram_107_tdata(m_axis_bram_107_tdata),
        .m_axis_bram_107_tready(m_axis_bram_107_tready),
        .ap_bram_107_addr0(ap_bram_oarg_107_addr0),
        .ap_bram_107_din0(ap_bram_oarg_107_din0),
        .ap_bram_107_dout0(ap_bram_oarg_107_dout0),
        .ap_bram_107_we0(ap_bram_oarg_107_we0),
        .ap_bram_107_en0(ap_bram_oarg_107_en0),
        .ap_bram_107_addr1(ap_bram_oarg_107_addr1),
        .ap_bram_107_din1(ap_bram_oarg_107_din1),
        .ap_bram_107_dout1(ap_bram_oarg_107_dout1),
        .ap_bram_107_we1(ap_bram_oarg_107_we1),
        .ap_bram_107_en1(ap_bram_oarg_107_en1),
        .m_axis_bram_108_tlast(m_axis_bram_108_tlast),
        .m_axis_bram_108_tvalid(m_axis_bram_108_tvalid),
        .m_axis_bram_108_tkeep(m_axis_bram_108_tkeep),
        .m_axis_bram_108_tstrb(m_axis_bram_108_tstrb),
        .m_axis_bram_108_tdata(m_axis_bram_108_tdata),
        .m_axis_bram_108_tready(m_axis_bram_108_tready),
        .ap_bram_108_addr0(ap_bram_oarg_108_addr0),
        .ap_bram_108_din0(ap_bram_oarg_108_din0),
        .ap_bram_108_dout0(ap_bram_oarg_108_dout0),
        .ap_bram_108_we0(ap_bram_oarg_108_we0),
        .ap_bram_108_en0(ap_bram_oarg_108_en0),
        .ap_bram_108_addr1(ap_bram_oarg_108_addr1),
        .ap_bram_108_din1(ap_bram_oarg_108_din1),
        .ap_bram_108_dout1(ap_bram_oarg_108_dout1),
        .ap_bram_108_we1(ap_bram_oarg_108_we1),
        .ap_bram_108_en1(ap_bram_oarg_108_en1),
        .m_axis_bram_109_tlast(m_axis_bram_109_tlast),
        .m_axis_bram_109_tvalid(m_axis_bram_109_tvalid),
        .m_axis_bram_109_tkeep(m_axis_bram_109_tkeep),
        .m_axis_bram_109_tstrb(m_axis_bram_109_tstrb),
        .m_axis_bram_109_tdata(m_axis_bram_109_tdata),
        .m_axis_bram_109_tready(m_axis_bram_109_tready),
        .ap_bram_109_addr0(ap_bram_oarg_109_addr0),
        .ap_bram_109_din0(ap_bram_oarg_109_din0),
        .ap_bram_109_dout0(ap_bram_oarg_109_dout0),
        .ap_bram_109_we0(ap_bram_oarg_109_we0),
        .ap_bram_109_en0(ap_bram_oarg_109_en0),
        .ap_bram_109_addr1(ap_bram_oarg_109_addr1),
        .ap_bram_109_din1(ap_bram_oarg_109_din1),
        .ap_bram_109_dout1(ap_bram_oarg_109_dout1),
        .ap_bram_109_we1(ap_bram_oarg_109_we1),
        .ap_bram_109_en1(ap_bram_oarg_109_en1),
        .m_axis_bram_110_tlast(m_axis_bram_110_tlast),
        .m_axis_bram_110_tvalid(m_axis_bram_110_tvalid),
        .m_axis_bram_110_tkeep(m_axis_bram_110_tkeep),
        .m_axis_bram_110_tstrb(m_axis_bram_110_tstrb),
        .m_axis_bram_110_tdata(m_axis_bram_110_tdata),
        .m_axis_bram_110_tready(m_axis_bram_110_tready),
        .ap_bram_110_addr0(ap_bram_oarg_110_addr0),
        .ap_bram_110_din0(ap_bram_oarg_110_din0),
        .ap_bram_110_dout0(ap_bram_oarg_110_dout0),
        .ap_bram_110_we0(ap_bram_oarg_110_we0),
        .ap_bram_110_en0(ap_bram_oarg_110_en0),
        .ap_bram_110_addr1(ap_bram_oarg_110_addr1),
        .ap_bram_110_din1(ap_bram_oarg_110_din1),
        .ap_bram_110_dout1(ap_bram_oarg_110_dout1),
        .ap_bram_110_we1(ap_bram_oarg_110_we1),
        .ap_bram_110_en1(ap_bram_oarg_110_en1),
        .m_axis_bram_111_tlast(m_axis_bram_111_tlast),
        .m_axis_bram_111_tvalid(m_axis_bram_111_tvalid),
        .m_axis_bram_111_tkeep(m_axis_bram_111_tkeep),
        .m_axis_bram_111_tstrb(m_axis_bram_111_tstrb),
        .m_axis_bram_111_tdata(m_axis_bram_111_tdata),
        .m_axis_bram_111_tready(m_axis_bram_111_tready),
        .ap_bram_111_addr0(ap_bram_oarg_111_addr0),
        .ap_bram_111_din0(ap_bram_oarg_111_din0),
        .ap_bram_111_dout0(ap_bram_oarg_111_dout0),
        .ap_bram_111_we0(ap_bram_oarg_111_we0),
        .ap_bram_111_en0(ap_bram_oarg_111_en0),
        .ap_bram_111_addr1(ap_bram_oarg_111_addr1),
        .ap_bram_111_din1(ap_bram_oarg_111_din1),
        .ap_bram_111_dout1(ap_bram_oarg_111_dout1),
        .ap_bram_111_we1(ap_bram_oarg_111_we1),
        .ap_bram_111_en1(ap_bram_oarg_111_en1),
        .m_axis_bram_112_tlast(m_axis_bram_112_tlast),
        .m_axis_bram_112_tvalid(m_axis_bram_112_tvalid),
        .m_axis_bram_112_tkeep(m_axis_bram_112_tkeep),
        .m_axis_bram_112_tstrb(m_axis_bram_112_tstrb),
        .m_axis_bram_112_tdata(m_axis_bram_112_tdata),
        .m_axis_bram_112_tready(m_axis_bram_112_tready),
        .ap_bram_112_addr0(ap_bram_oarg_112_addr0),
        .ap_bram_112_din0(ap_bram_oarg_112_din0),
        .ap_bram_112_dout0(ap_bram_oarg_112_dout0),
        .ap_bram_112_we0(ap_bram_oarg_112_we0),
        .ap_bram_112_en0(ap_bram_oarg_112_en0),
        .ap_bram_112_addr1(ap_bram_oarg_112_addr1),
        .ap_bram_112_din1(ap_bram_oarg_112_din1),
        .ap_bram_112_dout1(ap_bram_oarg_112_dout1),
        .ap_bram_112_we1(ap_bram_oarg_112_we1),
        .ap_bram_112_en1(ap_bram_oarg_112_en1),
        .m_axis_bram_113_tlast(m_axis_bram_113_tlast),
        .m_axis_bram_113_tvalid(m_axis_bram_113_tvalid),
        .m_axis_bram_113_tkeep(m_axis_bram_113_tkeep),
        .m_axis_bram_113_tstrb(m_axis_bram_113_tstrb),
        .m_axis_bram_113_tdata(m_axis_bram_113_tdata),
        .m_axis_bram_113_tready(m_axis_bram_113_tready),
        .ap_bram_113_addr0(ap_bram_oarg_113_addr0),
        .ap_bram_113_din0(ap_bram_oarg_113_din0),
        .ap_bram_113_dout0(ap_bram_oarg_113_dout0),
        .ap_bram_113_we0(ap_bram_oarg_113_we0),
        .ap_bram_113_en0(ap_bram_oarg_113_en0),
        .ap_bram_113_addr1(ap_bram_oarg_113_addr1),
        .ap_bram_113_din1(ap_bram_oarg_113_din1),
        .ap_bram_113_dout1(ap_bram_oarg_113_dout1),
        .ap_bram_113_we1(ap_bram_oarg_113_we1),
        .ap_bram_113_en1(ap_bram_oarg_113_en1),
        .m_axis_bram_114_tlast(m_axis_bram_114_tlast),
        .m_axis_bram_114_tvalid(m_axis_bram_114_tvalid),
        .m_axis_bram_114_tkeep(m_axis_bram_114_tkeep),
        .m_axis_bram_114_tstrb(m_axis_bram_114_tstrb),
        .m_axis_bram_114_tdata(m_axis_bram_114_tdata),
        .m_axis_bram_114_tready(m_axis_bram_114_tready),
        .ap_bram_114_addr0(ap_bram_oarg_114_addr0),
        .ap_bram_114_din0(ap_bram_oarg_114_din0),
        .ap_bram_114_dout0(ap_bram_oarg_114_dout0),
        .ap_bram_114_we0(ap_bram_oarg_114_we0),
        .ap_bram_114_en0(ap_bram_oarg_114_en0),
        .ap_bram_114_addr1(ap_bram_oarg_114_addr1),
        .ap_bram_114_din1(ap_bram_oarg_114_din1),
        .ap_bram_114_dout1(ap_bram_oarg_114_dout1),
        .ap_bram_114_we1(ap_bram_oarg_114_we1),
        .ap_bram_114_en1(ap_bram_oarg_114_en1),
        .m_axis_bram_115_tlast(m_axis_bram_115_tlast),
        .m_axis_bram_115_tvalid(m_axis_bram_115_tvalid),
        .m_axis_bram_115_tkeep(m_axis_bram_115_tkeep),
        .m_axis_bram_115_tstrb(m_axis_bram_115_tstrb),
        .m_axis_bram_115_tdata(m_axis_bram_115_tdata),
        .m_axis_bram_115_tready(m_axis_bram_115_tready),
        .ap_bram_115_addr0(ap_bram_oarg_115_addr0),
        .ap_bram_115_din0(ap_bram_oarg_115_din0),
        .ap_bram_115_dout0(ap_bram_oarg_115_dout0),
        .ap_bram_115_we0(ap_bram_oarg_115_we0),
        .ap_bram_115_en0(ap_bram_oarg_115_en0),
        .ap_bram_115_addr1(ap_bram_oarg_115_addr1),
        .ap_bram_115_din1(ap_bram_oarg_115_din1),
        .ap_bram_115_dout1(ap_bram_oarg_115_dout1),
        .ap_bram_115_we1(ap_bram_oarg_115_we1),
        .ap_bram_115_en1(ap_bram_oarg_115_en1),
        .m_axis_bram_116_tlast(m_axis_bram_116_tlast),
        .m_axis_bram_116_tvalid(m_axis_bram_116_tvalid),
        .m_axis_bram_116_tkeep(m_axis_bram_116_tkeep),
        .m_axis_bram_116_tstrb(m_axis_bram_116_tstrb),
        .m_axis_bram_116_tdata(m_axis_bram_116_tdata),
        .m_axis_bram_116_tready(m_axis_bram_116_tready),
        .ap_bram_116_addr0(ap_bram_oarg_116_addr0),
        .ap_bram_116_din0(ap_bram_oarg_116_din0),
        .ap_bram_116_dout0(ap_bram_oarg_116_dout0),
        .ap_bram_116_we0(ap_bram_oarg_116_we0),
        .ap_bram_116_en0(ap_bram_oarg_116_en0),
        .ap_bram_116_addr1(ap_bram_oarg_116_addr1),
        .ap_bram_116_din1(ap_bram_oarg_116_din1),
        .ap_bram_116_dout1(ap_bram_oarg_116_dout1),
        .ap_bram_116_we1(ap_bram_oarg_116_we1),
        .ap_bram_116_en1(ap_bram_oarg_116_en1),
        .m_axis_bram_117_tlast(m_axis_bram_117_tlast),
        .m_axis_bram_117_tvalid(m_axis_bram_117_tvalid),
        .m_axis_bram_117_tkeep(m_axis_bram_117_tkeep),
        .m_axis_bram_117_tstrb(m_axis_bram_117_tstrb),
        .m_axis_bram_117_tdata(m_axis_bram_117_tdata),
        .m_axis_bram_117_tready(m_axis_bram_117_tready),
        .ap_bram_117_addr0(ap_bram_oarg_117_addr0),
        .ap_bram_117_din0(ap_bram_oarg_117_din0),
        .ap_bram_117_dout0(ap_bram_oarg_117_dout0),
        .ap_bram_117_we0(ap_bram_oarg_117_we0),
        .ap_bram_117_en0(ap_bram_oarg_117_en0),
        .ap_bram_117_addr1(ap_bram_oarg_117_addr1),
        .ap_bram_117_din1(ap_bram_oarg_117_din1),
        .ap_bram_117_dout1(ap_bram_oarg_117_dout1),
        .ap_bram_117_we1(ap_bram_oarg_117_we1),
        .ap_bram_117_en1(ap_bram_oarg_117_en1),
        .m_axis_bram_118_tlast(m_axis_bram_118_tlast),
        .m_axis_bram_118_tvalid(m_axis_bram_118_tvalid),
        .m_axis_bram_118_tkeep(m_axis_bram_118_tkeep),
        .m_axis_bram_118_tstrb(m_axis_bram_118_tstrb),
        .m_axis_bram_118_tdata(m_axis_bram_118_tdata),
        .m_axis_bram_118_tready(m_axis_bram_118_tready),
        .ap_bram_118_addr0(ap_bram_oarg_118_addr0),
        .ap_bram_118_din0(ap_bram_oarg_118_din0),
        .ap_bram_118_dout0(ap_bram_oarg_118_dout0),
        .ap_bram_118_we0(ap_bram_oarg_118_we0),
        .ap_bram_118_en0(ap_bram_oarg_118_en0),
        .ap_bram_118_addr1(ap_bram_oarg_118_addr1),
        .ap_bram_118_din1(ap_bram_oarg_118_din1),
        .ap_bram_118_dout1(ap_bram_oarg_118_dout1),
        .ap_bram_118_we1(ap_bram_oarg_118_we1),
        .ap_bram_118_en1(ap_bram_oarg_118_en1),
        .m_axis_bram_119_tlast(m_axis_bram_119_tlast),
        .m_axis_bram_119_tvalid(m_axis_bram_119_tvalid),
        .m_axis_bram_119_tkeep(m_axis_bram_119_tkeep),
        .m_axis_bram_119_tstrb(m_axis_bram_119_tstrb),
        .m_axis_bram_119_tdata(m_axis_bram_119_tdata),
        .m_axis_bram_119_tready(m_axis_bram_119_tready),
        .ap_bram_119_addr0(ap_bram_oarg_119_addr0),
        .ap_bram_119_din0(ap_bram_oarg_119_din0),
        .ap_bram_119_dout0(ap_bram_oarg_119_dout0),
        .ap_bram_119_we0(ap_bram_oarg_119_we0),
        .ap_bram_119_en0(ap_bram_oarg_119_en0),
        .ap_bram_119_addr1(ap_bram_oarg_119_addr1),
        .ap_bram_119_din1(ap_bram_oarg_119_din1),
        .ap_bram_119_dout1(ap_bram_oarg_119_dout1),
        .ap_bram_119_we1(ap_bram_oarg_119_we1),
        .ap_bram_119_en1(ap_bram_oarg_119_en1),
        .m_axis_bram_120_tlast(m_axis_bram_120_tlast),
        .m_axis_bram_120_tvalid(m_axis_bram_120_tvalid),
        .m_axis_bram_120_tkeep(m_axis_bram_120_tkeep),
        .m_axis_bram_120_tstrb(m_axis_bram_120_tstrb),
        .m_axis_bram_120_tdata(m_axis_bram_120_tdata),
        .m_axis_bram_120_tready(m_axis_bram_120_tready),
        .ap_bram_120_addr0(ap_bram_oarg_120_addr0),
        .ap_bram_120_din0(ap_bram_oarg_120_din0),
        .ap_bram_120_dout0(ap_bram_oarg_120_dout0),
        .ap_bram_120_we0(ap_bram_oarg_120_we0),
        .ap_bram_120_en0(ap_bram_oarg_120_en0),
        .ap_bram_120_addr1(ap_bram_oarg_120_addr1),
        .ap_bram_120_din1(ap_bram_oarg_120_din1),
        .ap_bram_120_dout1(ap_bram_oarg_120_dout1),
        .ap_bram_120_we1(ap_bram_oarg_120_we1),
        .ap_bram_120_en1(ap_bram_oarg_120_en1),
        .m_axis_bram_121_tlast(m_axis_bram_121_tlast),
        .m_axis_bram_121_tvalid(m_axis_bram_121_tvalid),
        .m_axis_bram_121_tkeep(m_axis_bram_121_tkeep),
        .m_axis_bram_121_tstrb(m_axis_bram_121_tstrb),
        .m_axis_bram_121_tdata(m_axis_bram_121_tdata),
        .m_axis_bram_121_tready(m_axis_bram_121_tready),
        .ap_bram_121_addr0(ap_bram_oarg_121_addr0),
        .ap_bram_121_din0(ap_bram_oarg_121_din0),
        .ap_bram_121_dout0(ap_bram_oarg_121_dout0),
        .ap_bram_121_we0(ap_bram_oarg_121_we0),
        .ap_bram_121_en0(ap_bram_oarg_121_en0),
        .ap_bram_121_addr1(ap_bram_oarg_121_addr1),
        .ap_bram_121_din1(ap_bram_oarg_121_din1),
        .ap_bram_121_dout1(ap_bram_oarg_121_dout1),
        .ap_bram_121_we1(ap_bram_oarg_121_we1),
        .ap_bram_121_en1(ap_bram_oarg_121_en1),
        .m_axis_bram_122_tlast(m_axis_bram_122_tlast),
        .m_axis_bram_122_tvalid(m_axis_bram_122_tvalid),
        .m_axis_bram_122_tkeep(m_axis_bram_122_tkeep),
        .m_axis_bram_122_tstrb(m_axis_bram_122_tstrb),
        .m_axis_bram_122_tdata(m_axis_bram_122_tdata),
        .m_axis_bram_122_tready(m_axis_bram_122_tready),
        .ap_bram_122_addr0(ap_bram_oarg_122_addr0),
        .ap_bram_122_din0(ap_bram_oarg_122_din0),
        .ap_bram_122_dout0(ap_bram_oarg_122_dout0),
        .ap_bram_122_we0(ap_bram_oarg_122_we0),
        .ap_bram_122_en0(ap_bram_oarg_122_en0),
        .ap_bram_122_addr1(ap_bram_oarg_122_addr1),
        .ap_bram_122_din1(ap_bram_oarg_122_din1),
        .ap_bram_122_dout1(ap_bram_oarg_122_dout1),
        .ap_bram_122_we1(ap_bram_oarg_122_we1),
        .ap_bram_122_en1(ap_bram_oarg_122_en1),
        .m_axis_bram_123_tlast(m_axis_bram_123_tlast),
        .m_axis_bram_123_tvalid(m_axis_bram_123_tvalid),
        .m_axis_bram_123_tkeep(m_axis_bram_123_tkeep),
        .m_axis_bram_123_tstrb(m_axis_bram_123_tstrb),
        .m_axis_bram_123_tdata(m_axis_bram_123_tdata),
        .m_axis_bram_123_tready(m_axis_bram_123_tready),
        .ap_bram_123_addr0(ap_bram_oarg_123_addr0),
        .ap_bram_123_din0(ap_bram_oarg_123_din0),
        .ap_bram_123_dout0(ap_bram_oarg_123_dout0),
        .ap_bram_123_we0(ap_bram_oarg_123_we0),
        .ap_bram_123_en0(ap_bram_oarg_123_en0),
        .ap_bram_123_addr1(ap_bram_oarg_123_addr1),
        .ap_bram_123_din1(ap_bram_oarg_123_din1),
        .ap_bram_123_dout1(ap_bram_oarg_123_dout1),
        .ap_bram_123_we1(ap_bram_oarg_123_we1),
        .ap_bram_123_en1(ap_bram_oarg_123_en1),
        .m_axis_bram_124_tlast(m_axis_bram_124_tlast),
        .m_axis_bram_124_tvalid(m_axis_bram_124_tvalid),
        .m_axis_bram_124_tkeep(m_axis_bram_124_tkeep),
        .m_axis_bram_124_tstrb(m_axis_bram_124_tstrb),
        .m_axis_bram_124_tdata(m_axis_bram_124_tdata),
        .m_axis_bram_124_tready(m_axis_bram_124_tready),
        .ap_bram_124_addr0(ap_bram_oarg_124_addr0),
        .ap_bram_124_din0(ap_bram_oarg_124_din0),
        .ap_bram_124_dout0(ap_bram_oarg_124_dout0),
        .ap_bram_124_we0(ap_bram_oarg_124_we0),
        .ap_bram_124_en0(ap_bram_oarg_124_en0),
        .ap_bram_124_addr1(ap_bram_oarg_124_addr1),
        .ap_bram_124_din1(ap_bram_oarg_124_din1),
        .ap_bram_124_dout1(ap_bram_oarg_124_dout1),
        .ap_bram_124_we1(ap_bram_oarg_124_we1),
        .ap_bram_124_en1(ap_bram_oarg_124_en1),
        .m_axis_bram_125_tlast(m_axis_bram_125_tlast),
        .m_axis_bram_125_tvalid(m_axis_bram_125_tvalid),
        .m_axis_bram_125_tkeep(m_axis_bram_125_tkeep),
        .m_axis_bram_125_tstrb(m_axis_bram_125_tstrb),
        .m_axis_bram_125_tdata(m_axis_bram_125_tdata),
        .m_axis_bram_125_tready(m_axis_bram_125_tready),
        .ap_bram_125_addr0(ap_bram_oarg_125_addr0),
        .ap_bram_125_din0(ap_bram_oarg_125_din0),
        .ap_bram_125_dout0(ap_bram_oarg_125_dout0),
        .ap_bram_125_we0(ap_bram_oarg_125_we0),
        .ap_bram_125_en0(ap_bram_oarg_125_en0),
        .ap_bram_125_addr1(ap_bram_oarg_125_addr1),
        .ap_bram_125_din1(ap_bram_oarg_125_din1),
        .ap_bram_125_dout1(ap_bram_oarg_125_dout1),
        .ap_bram_125_we1(ap_bram_oarg_125_we1),
        .ap_bram_125_en1(ap_bram_oarg_125_en1),
        .m_axis_bram_126_tlast(m_axis_bram_126_tlast),
        .m_axis_bram_126_tvalid(m_axis_bram_126_tvalid),
        .m_axis_bram_126_tkeep(m_axis_bram_126_tkeep),
        .m_axis_bram_126_tstrb(m_axis_bram_126_tstrb),
        .m_axis_bram_126_tdata(m_axis_bram_126_tdata),
        .m_axis_bram_126_tready(m_axis_bram_126_tready),
        .ap_bram_126_addr0(ap_bram_oarg_126_addr0),
        .ap_bram_126_din0(ap_bram_oarg_126_din0),
        .ap_bram_126_dout0(ap_bram_oarg_126_dout0),
        .ap_bram_126_we0(ap_bram_oarg_126_we0),
        .ap_bram_126_en0(ap_bram_oarg_126_en0),
        .ap_bram_126_addr1(ap_bram_oarg_126_addr1),
        .ap_bram_126_din1(ap_bram_oarg_126_din1),
        .ap_bram_126_dout1(ap_bram_oarg_126_dout1),
        .ap_bram_126_we1(ap_bram_oarg_126_we1),
        .ap_bram_126_en1(ap_bram_oarg_126_en1),
        .m_axis_bram_127_tlast(m_axis_bram_127_tlast),
        .m_axis_bram_127_tvalid(m_axis_bram_127_tvalid),
        .m_axis_bram_127_tkeep(m_axis_bram_127_tkeep),
        .m_axis_bram_127_tstrb(m_axis_bram_127_tstrb),
        .m_axis_bram_127_tdata(m_axis_bram_127_tdata),
        .m_axis_bram_127_tready(m_axis_bram_127_tready),
        .ap_bram_127_addr0(ap_bram_oarg_127_addr0),
        .ap_bram_127_din0(ap_bram_oarg_127_din0),
        .ap_bram_127_dout0(ap_bram_oarg_127_dout0),
        .ap_bram_127_we0(ap_bram_oarg_127_we0),
        .ap_bram_127_en0(ap_bram_oarg_127_en0),
        .ap_bram_127_addr1(ap_bram_oarg_127_addr1),
        .ap_bram_127_din1(ap_bram_oarg_127_din1),
        .ap_bram_127_dout1(ap_bram_oarg_127_dout1),
        .ap_bram_127_we1(ap_bram_oarg_127_we1),
        .ap_bram_127_en1(ap_bram_oarg_127_en1)
    );

endmodule
